`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mWsTIr0hDumHIrVL4Sph3sZnrExdfvYUaHHEQ+XvKp3WoEMgbuc8wI6WGdF+aZXd74dP0VU8CDJF
rTc4wjr8og==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TxaMRpwVT3dY6PSvNCGyS/ahlYjOrJJmKT+BNylJN5hugjKGMC8/1qXAVVGRpwV2FuSA2Pklc3fT
WQbShwV0rCE+dPsF79sOHd/1f/A9IleIhJDOzcJzz+3mL1ioxSXyoZUBEGTecDW8nc3N3+B65SkS
DKBmMACGu7/mINFoNHE=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JC8mAxsIlFRJGmj17DZdjH4mH/Vcs9yPb0kKkuWCYAHCr0wQsgeL4wCtpCHyQbGuWZ+PBEP9JhhX
rgGbU2uJf5GLE5fIAJX2cjVEdSxgICyMUKBn9iWJ4qA+Wr4+NSIRsYXyNG/klviSkYFj8R8xqBi4
JIU0it7GFd5owzw/N48QrTtH9JPxqaWOKD0Sz7xYgZupHbU9lz2wQ0AQNICLysNhpo9wXGByQVPq
0lp1SkTtMO8yFWwBadKsOH0TEr4CnrcA/eYRTci8MzIp6geTPkjQrPd1tCgKMstoBnSlPvs5Y2ST
Sduv4VO+dNeOL6ATNzXdaOlAA3+N1Z5Clakjug==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gKvljGb5SdLpiA6Eldy+lpgJczSDlWQF0b9oTmyxNzAildWi6WTIuzPRDD5g4PLoGt2ze4j8avF7
A3rlK3R3I/usUDtAlXhrJVq/QheQ8PqmpWge4Xk26cl4/zBXCjg19Se6zXRyLGfJJY2oH/+O96kp
2FJTXdXUeMl4dR95s5R1VCF7pO4NRwt1nQ2XvIr0UeIuz8X2X/sycix3WJ0uCmKfUFmL6SH5coQE
BOqjQG9cWwje1BjNAt/sAYzFB7089h7l8VQxumhnec8rLFnvUl+UgZPl6DsxgojlkXZsJH9Zks+4
9WCLstyjUTxYupGfWmM4QJOBeEg8y7bKui2OOw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kYioazr5SJAGhsfiAYbuRNcRbGN1OtzgOrMIZs+TO58HdjgS4YuQQUw0OnQJobWLk+Md+uLUyEcg
y9+zClYvGXkMWvOoFMKD9la+NfcWlcx+UQhM/zKI+fK2HoYAUAMuMyqzC/O3UgqkiFaCnCzQgFKl
RoCXLHYNciLdax9PfS2K8pHyecwcRQPbKHXqdlpnX6TIwRA+rnhK1mKwWKoqBni4mLhsCYkZ7UUF
f5hEfcyQg0asEhmXuVLv9Xa16TQ5DuUvXi5Mv/9WhXvcgtT6HMN+D/WSwvDzkG+QmJy2IRSBGlOU
KQEAGtoQuBhfYuD23aoTAJ7ZOQsVGG/SwEINhA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
utn/12CyyOQ44wwHDcCSmCaG3jtXJ3Ca/LQ1iendDcWJxAU0Eotu1FV9hECpT6yGaMqQkt6iT4gn
po0qm9CSYNuxlJ2Y30iOIf+3K0KttEZMcba6/vg9u8M80bH9rPfT5HKG7g5A7+DpIWBW+z9rl5px
g/6m6ofDqoZiS7OV+YU=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qIs9eGqa1hcoEUiz8xnByjZfZrMrFCy0vpL19y69gHwBwXKHLzswY/tTb/neH9Dl1M/yKT+UyxVS
1Wh26oD6KhUsHxJME6BIovM75ch4lWnRb20D5AWZBTRxTt5dyMAiUKWAepHP4z7l5XGfKxHejYLr
vPvIG/gCeO1XlcZhZoOIy5JDZSHu4clHstIbsVWzWZeAbP/JtUDBV9HQyIGL0u/a6HCatIFUsbjh
A7C0YQ03sLaa6Y4Iu4L6I4sVltdxiPCGToQVoJOyPG7k0xRCIP2HCOPZprQUP8b0nBUuGWqh8I6j
40Bpve17+XnmaaZCeJcru9qtndakspqS56Hssg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 98368)
`protect data_block
PCxoVWOuPJAoh2svws1LdI6h49LzgTd3Emybc5SHzE+Avq0vHQ0sHsjqiq/XasU4Bv/bZa3u7hhZ
S9ymexJqVHoVWqoLGGgxzBfP04m1gFAqHpD9CT0y57H4VrxCPUZgHIIZmeGCFMvCnESFHBCwk5Ku
KEIrI+5c8TeqDMbj+pKrG2MnnKfQ12z+WGycH+a0snG/ZnAUlzxpZgymA9gjx1XBaBMKU2NJTcmU
Qr6AffiyFt1YUUftAgLuh7PLtR0ab0hpDTKgY/MtGbFlLBvnAs4mmyfAfRApl8eNGpzF2UUkpkSt
OgHUsIE+zvg3BEu8OqG3xPY1avUz4+lHzwwXeoEWLrV8jN0gwdIBZCsyePKpmFWxYgPE/tVZg06W
Doe4/3r1AnjziGtjc74OpE2sxyIzhGIp2n4yMVB1o3lorigtb2llecnhF4VhVZAbecElHFmbhhJc
ebNx8SB220Y82aRrMF9SQTkmz/Av5w17BIv6xnvmz2B2IOgcfYx5yxdfEHDlwcBNQOHnINOmfcUd
rXp/T0QgevmayG0PtqcB8HEU61bHc06QIU/FSxy2BB/NgsOyx28sJGnIO4eEpattondcPyVzqr2E
zGUollenCZmBCy+W+aRjUAjtvZURCDh/adjvadeiN8ycMB73IP2xzy8/emE1Euccilc+zzoWILUT
8YcaC2846wMQ4PM4SNBcaF2AjEulbimwHPEroPAz3Qz0qvzM1SAO42TJUFh6YytGrp0CRFzMCJHn
CXxB1UqsVEcbWO4clJPT15rVTXrGoBHXCicRJfEMtkBcirNzCi1kRH9B2nZ0p6xRPeYK6i97pUK4
D3dxgJ6QSbFdlCVvbj9pluY0UwBNydCTdVFm3325I57UDpffYScT8WXAh/6zGGs0Jrk1O1m8TYXM
W971BourEUsKwk+QTTCPhMt03cYKFfRbPDAcLVR9rnKoD76MDXGxUtT1l9rLf2iqFQAMTWgFRcCl
L7i+joKLvO0tnuVVUu6c96SNI+sslEQDnOTh8iVaReUDHzz2TLFZS+cAfbhN6tf/FBqwJUVd9Af+
51BWc+kd4EO1FKu38l5vRqmEScr6G4ApQn+J5tW6ut4NvPrSI5fM29IOhPNkcD2XW9hEZyuXoO9c
if2+8goIXF44Sc3r2KBXI92AN8a8KOptEJarxEQfx1tt5VyalN7dKY6I57cpUwnAQQdyuJstS0BG
JE1HIZXjBRYLG/tHPhiBpsM2pd8uvn/vKjb2kUhV/7Wgi1NP9IfvPp2mWDUNlnogBcrrol+qOtVE
SW63MbNZlHh98eny4Du0Qr4nFSGSlk8r/Z19EwohI2pRONOPNhOhsIajyShk89vbHLdX4X15shJd
bPb3slQ8jeV6oJkQLzAA/ocLNBk5dB3e01U7FIjhQ36JgxCdeOcJMwFfzTTUx8ftG1fZv0yxpvTb
XAauOWHt0Rdoufrx9ESAowQAFtaoXcUwunKSmsopPWHfhQg66dfUaqWRs7OiIfodrWdbV+dp1ImY
2Aft40yqcUoNSNJ6/sUeC7q0lgJY24XSuocVLem1hpT16b7pl8I3cLtnTeQ064TV5rP6DUVIcz4M
FCmuuZM1LOYL+qEpUxO9pZIYaD9dOFZgjRI7N/h/UykQXE45b0KShGl425EY2eF6CLgmiy7h+b/M
UHrPz3yOMV+EORuze3i41cjV7rwERGU4wBScUUkuRcOAY/LUh5/FuNwD7G8sCXFyey9DFjjWHqtQ
RPLJi/bCeZoE+HTfSdxtePRgeWW17TjCRyufX1wNHfgUVre1ut238SazwZSgbUsxylb/UUGNDRlt
Pw3kcZkvwOAPOWeC9gxBKcsFeXT5yG3x2fMw8V6zt54JgbGxhd8RobOBkPfUyDMCPCgER3tzILAy
gos03i5pnLIa3BosnSLBkY+TKd3eo29qqiRqao5mHdeLoZSlnznXXXZnKiKX9Vz6TvEj3C+YqEA8
Pn4ttKlsRF8fseRqvY7ICgmtH3EjoIw5apb+AE5H743ySc5szVtuf+2hQlNj4FmTe9Z+t9wSxm5W
L5j5jpvFodWjzsSPv4/9yPQD0yVRPjTZ/62aJKZgYbct1Ki3+mMhs9Om3soPwik1rFaFhFEzi+o6
daWw+uxnWlrTjcALMTGO5OES2HKY/Dtmwctxyy3z7E/6FzPvSuSDruBCGDG2RY09QdqSg0WEMhYq
pJ5CvsKShPOYGs/ZPLoz6y8U2F5z80QbkjVpqxMZXRFdseW9PbjwZ5IjB8J5bYU10qSE+A1fY132
PqEOs505+rg8jNe6y/sx4oxcSDkP3q4rH0hfJWkrCgOv8GVKk1iME8cog4Ri8oeZoBoxdjctDZSI
xD4tYEVS7wTI0fyHVgRDGrBHMP+LmyvzT1Yu6bNE0eiMtI6WzDSQ8/8nt2PliFC17m4dZX/YGXtz
gtiQfysj+od152hvfTRKvfssJQqpnvzpqajhiXngwakAnsxYjrxx2S12PBpCzAW3m0VbrVC8cgOD
27oScW7ILEq0QIS1zTd84XOEWmdCW1+lBWHhTaP/sHnw7dKS8pmt/kjzSrakBsBN5ePL57PWSLSg
/zma71qzXawQ5JxZGV2cpPlHTMAKoyQOhsJws1Jlti9onLc1pzx55ZQHL0nlHr8SicJ0lq+v5Ic7
vY593Lmwnr/XQwnWtB2KWs9aXNSxM1Opw0kdTrQXwlVb2RWfHp2R80YxZIz4uA5C7L6qQi3PRDej
wYL9kjZpKdulAX3yJHQrqqWspFb4n8N3qaWTDMJiluB2YHxrSgH7oOC8iCV/euriWjd9r7BBszou
rq3R00TM4r7yYeZ5554n4eG/NWO7aQhVrYy9eTdsqF7VWjUyc5kSCcIi2fo+hvcj9337uMVwoQUa
FhD/ZVNirJJWbQOp0LnLJS8TSWFwWqt4jVTItdYFt5O4Tw66r5ZYW2bJ8K/wh3SWbCEy/9LSYF0H
vdWgdzKvMHUERqyqxyl5ViaAfagUWXYdlJFb3oyg0bEAbgqlRBVRo6FC12IU0Ihu5nKcI2VxGM1m
nZ4bvOp3Y1GdO1nHePNOFBpMdOlzbmLuiuMhy0gzCIQWRiv0Iexig+/qZCxLckakV4qLz4lDZ+pH
fItQEp6XnOYb6GZiEm7kKtNimA+acmudsIfzdMLdssIIyG9lUzprxWQr60UCIAWapp1Ne2fbrCg+
JAWKtw35zz3QoZD1E+BscPQTrggj2JdIZ+LDmVxebTlGCJmmIlAE/99pTzQegPiCUCZmFP04/5/a
QamX5OgfLk8Shx0aSp7Nkj+mq7Kd8mbXq/08BKz8+DzxZCeMFDU9AKelxzk10HZ9oKalXDPkH0Gp
KUj7trFlkRd4ubpwqb9/pO7ezMihDRmQsLbRGP7ufiOEjjbG6jqFGsLPez/1dfpqcV9ITejI+Ugc
gnKiRUqKX4OG7tych8lzCsAsKN6ztin2gK7PocUeET8sxGsBJUcOYwWzM6eOVfncI2xCBC6joEby
/WazGTNcxfGa9r3+lDG+EXIiiZ+dAN2LjfYLKSXz57FL/5PfGONmoKzv99+eHaND4MtKx06LBHNa
XK9ekn6D0VIFBgzscLa/nAiVL8MCZ2CWKNhIEB5U4Lcdz1kQIqMz74kPhnNcS95UQeGvHI3LWHoy
naEP4PsmYT4JCT38yJsZ4iEyZErmzIzEwzzebz0GW+6hh0Pv70ulFPQbj+00fgDr32jm4XiMs5yF
vSDhtbhhOTeyXrbo2xK1lkKWpi+PZOxAbkXGdOb/cgop6LjB5Za5ZUdSPfrgCmy1SU4yMA7Ev3gK
a9DLOB1dljazi05NWCsOm5Tr3DVbhl00fMEiWbG+/qNHfWVj53cU5Nmv+qqoMGKBj25jDUieuGt2
vOyPYTQn0uxJeE+czhaKgrlYQWc9pUtGeadYVr463Eia8JPLwB1Zf7+GBnwhjHM6y1noAz3E9iNV
gWpVPkZTXU9oGtRqn9XuFAncjVbwb+6CJCFpLx5OQTVotNMw4ewMeUxp7UImRyeHfQ0AP7GmgL/3
Z7FJ13V5GKkg2/V6tWL8pccjAjOH8prFyHY9WRS4171t9vhau95BwDy5z/n/kAHJTczqeuycKqMW
jEmKJVcefwjp07cuQjpubPl+0m8cqfUbyuJBWJ+mUzPM6nyF7tj9lrzPB1EYVMK5e2Q707Ws4+KL
15rZA5JAYkWa9t0JLU42VvjQrspuBzFdHM/I0P109ZMawsly1GQrDJLs6vSeoii5INZwjBBgi6dp
NvANZ9oxBkiw/dm2+FJXqeyukrLNljMW99Gijvkyvfl0BM7wOjqC652TstKWbpTEIoRdv5WCzHKR
IiOHu7EG2InBsP4G1ye/LVkxSN1EJ6xh0HYGbp8Pu1KTRvEgc8HrgYDBGJE5amOluT7/v2/0B7es
FgyqYli8b2jTN+jd8N7Ka4Z5cPTpcUME9BpnYPP2wu+Yw6URDSF9kRpIclaRv56AXXzBKVtRVKU+
Dyidzct2f4HOtvaP2FHRaYcdVY9Z9Nn1pG8Y+GCXYqqkPsnYDBpTC7MHLQcV8Jb8glPfLKX57j2y
mxPgXMrQ4Yf64cCDrDNUw9G3lUlqrrmPqmJTflGnVAQln92YP/S4YqIUAPNvePomBkx/5/I5S7zF
/46hRB69/WgloboyyV5NGp7F87x8be8pnu0/sQuEjV4t4aSGyuJocBLBsbV8v/tV6ADz6BcoEGUQ
5/FNKHsDBUewjytWeh1a2N0GtVrWAKjaNxls1VpygwqMt7mSZorhNPhQjY93tsfYFzguGppDEKC7
aCWqUf/kku8UW3EyOngIW9b7L3578dBcRV5+runkiTvYL6jwzn8ExuPIdE0LnHm41pmQbirBJkvf
mQlJNuo9CmnxE/8IeZhtft60KCokYx+Iss6MBPJb2Q/BtvP+/HG+KN31bd4uREoaeUrifogtk4iB
yNKvisSKl0KzGxAycGlzRUcQyxqrDhO6aO+3W58IMdHUBDEoxzPfPrIy62FI5LuRUYphz99pp1Z/
iCqqA1HLPNTOWJA3/t6JgHpcyKAnR6dDbAY5zdi1KSUGWqscA0f1pvklPJGHOMjWNaZQJBEmNqID
0V3Ztp8oIYfMDxUUiU1NaQodPz6iCisH4ZJSCFIwJh6/F5wu0WMNkfEuRmhvpFULr/pkw3h4dGdW
4r65LAOSJmy7L0BBd1GTJqcGsIzOlflmRM5WCsZ9NfXTxZgeCDFxm/RNcNX7QWcEOtTJjCBr2D0u
S9u0yE/KUIOO1yFQyFXypb/ImUQA8++51xtjmlNh4Wq+t08nud5CcPqHav1x9Nu0DPvkKG7++m1S
MWcKVnD4vCHSv/37Nw+nVJ7o4LNmmN5imtHuJCHBiKryjU+eNl5H4nrqkhApNMtXdm20zGbsMjvv
5xOWRmHtS+7AUTYH8rLzl11YoZwdEshzTdxMS9j4bdSlISa8aBDvwxM3/HIwIaTlI1WbhvK91KlD
H82j3HtgjPx8pxOI63nmjfBjgvr6tyLOfY5tC9w/UhksAlvGcMcdxqAsTEJzFqksQhzji50vriFl
GBMB+Pgu1wLqaaRLx7nY5CCmsO2/7RvamDxhns0emIGWxhzjOap6OV1r3uUg8EtuU4spJV+7svtp
RDdilj2Bsly2RMuWESPOrkUMJfW3k3csFbPB94W3VdSXyZrhdZ9XqhYNcDHanO5Wglu78Zw2lfcB
uP0l97X2qiMjFl/n/wrBSPA0v1TEoXOdQKxHVTy+8/r2XhdGkaDWQeMAAEnky9jCYHVMqa66IJjy
Oxlx5mi1kXyjZFeS+xGWtc6K/JcxBMM2ohEog3k1zf63KgOTdBN0AANX2JPhrg/P+MkugTNd2klG
M4fR8tThqsICYuKCt/7i1jl9zEyj5coR4hk+fW+IqjyOlggc5qAUo8uZkaSJt7moNBS1VRDUXXFe
StM7cgekOV3Yp/XHJwBL0/YYlTrgN6MAFL1vRHZMExcGuShyXEC2oNwaJSnTHhkSt81Zzmj+Bt7O
19YS4khduyS/J700VTY4tbXLyOy362QYqu5UCl09yx1TEZKztYDlBY31CJV2VPtMIxpQPsAKtz7p
vZgXIE6KgL5x5dSVpo/lnfDCjOsiiVUD2ovyGNbwO/YULlaRyUoSB+kA+4Su2JbRT9SoslTnVXg6
6tuySqv+XvSywky4oKY1JsFCo1ouBv8EGBkA79MgFzu8XFa06XptWo+AapX8UTojpDv1xYgIxmdD
GwaW6bGIzLZYYrkvD9ot3Cxvjcm7k9lgVjeHFkT0btcbEGVJPf4ykPvGxQkUiCWufJ202Xjn3I2O
3XSTHr5OtTa0h7GVIzUYA636AlzocDICtgKTiM1k5XDNT08TUK8FiXp69O+xImBVu8YV1INL76F6
HHJF0wclWD835ja5Ub8TdVuU3zX7denlB6tfGGUlAj113uskN4jbtn7KkjpRKgB0xaBFQIg5HgUV
G9aKbVDj6JLYGUOz839b3WdGu/Y9diKUtoPWk3ZviM/QkTnJYjoOMQvGPUHhyf7H5EeHWrs75A5n
vljsBjgzuRHHU1IlyC5ScOcqxRPqODJWtvPh8Z208wfp7VTamkkm7C1SajXXv+yVoMFLFeYCi7eo
GBYynCddNjHSu+vdbmRpVyQjO9vEbxRGK8yPoC0T9rmuI+KYK9sEH+VsOcxcaP7AWdWLAtPHNsI/
MVO3j3WE+hNNR9UnMJwehpmlCfKRs6lR1YDEeX5rxhefK297SGfXkAvaOVeidCzb6pjM55e3GeNe
PQ6zsrvr2K+257gKpaff/rJbshUO5EEF+HwF7+uKzg7CmcivZz3JMj8BN7olIGOkjmBMaycIqU4D
MxoVg6ns5Y5jTHcHBgMOZ7gTNaKmUJqQrDUTadNDtROWQ4p6rwLazSOayxEGkWWY3CasrnqdAGpL
rVnKKfBHtoWv6X5Q6lqCe7aApKEVpDm5ljr48i9gdF3tGLMyT+adQ5feSNhMAorGUWWxSS2WVyCI
2w/ldqavfbwVXyLNN2WIbpifEyBCRCJ60LydFQPSlAzZX511MV+oO4zfOAEdedCAxpYQ71xjf0v1
a5ORByjIBd9MAlClKV71aRwaAdSp57o7NQft8adX78UO8qvRTZaDHOSzMGvU5BqVTtEwl0hG8K9K
gX6bM3jIWutTigI9w6bQ0wHF4GlbYgIN4IgL+JxuaeCt4VyqDCx3EUHKzfu32zUvFY1mRQzhG4Mu
T4wPRy1p54huAy9diMZULeA7oEq8OwcGU/sIKP9G3J27FKZM/IFAIuTD/IqnPbBD+qZJ6RgXXq4l
q2HHfVUmrksFWrOsWOhCZfqI83sPrP3d3UpTO6LknmpqjkbPpiCA8xZDJOsO3g/VIVk1PfAugHVL
6/aE+ffUmreX6IGnZWOuMnuWr5M4s2ZcsT+VVQVgzBmrIjLFfkjrXykFEbqCjq51b3W4bkGR2Kgf
FrGbxpyRjALJPFdDbGj1G+yafBS+C2UREN08JYNnajjEd5tumsPPBYzlqNZwagcaYKyuHsMrpB1w
nsDyaMh+PCsWat96zTQOqUWhmEDmd5gq/FBgMc9BDtqqGW0OA0Zp/0L22Psc9ahToasfSBR//LSD
mCQXBprIj/zBOPPr534Bi0fcxUWKEkY94eS6fZ/WgflvohsM2/TtpFqCoXDwymXnAO8z5REOohYG
soUzupuVo8HHb9EtrnBZuWehNO4NJsKMuEueHVDK0DYSfZz6lbn4Za6wiMKe9TB6iwwL5ySse0ny
ZP8sgd5OiFEP09pYrFP67+HH9V0v8TQ1ALaxhtXw+fnTAVs9V33uWuN6vmVmn6YNFr3luKuzbsIi
C5pYyoHtAwUyRV6I4inAHQrN4PWzlP6wu1ZNz3uSjhfmNHI23z02VK4fyWnhCZ1t15l/8cGfj53z
xULlKvyU+4G+jwB72QnbZDe57NBFqK8Jm/S4guGaLYX7ZTTVYVBryNPl8c7gbny9XpcKkLVdwbk1
Sb8+nLK922GVCQzwMWSZJrHNZN9Xj6y976cwL4l98w2cykQ/HC7sUUJIdJNisn2uMVBZSYLa6ZJ+
/G2Shv+R/WxJFba+GGbl5yC30qXTu2Vl34Zum0IDZBw/VOXSHaG903sxAsBRay7CCAq//7KTkC+5
JaLeK6mx5e1BbN7MBnbgIM2i5NPSLhpRbZYPCWHGdzfdiLBzbnz0MFVJCOJzL9AehtyteWNJg/Z+
up60LHuxpNEJi13cpOdlB9lvHJQCnFtg0V2RMQ/8SM6z+gen7ZftzbbIE3koWPdZaiWFUwcBA3V1
eD+AviLOY1SZItXvJ4tdnomYQBWDJLZQRuTg3ZCZq3aDytysm+he6sLrJS1+o0hDn9d1nm0PUJ2x
NX73fOg3NT98vnGHSLAeN6XePqvZwkgSULz5oWF8hwxjB1p6dh5GakVfJQOY6961+Wep4tEv7S3c
HZWkF0jA+VDI7XGZnCsepjZ7z1j/AWu0WepTHi/K93s3vkhqL/T7ryUzmPUomhtc/HrKocbyRAGI
fahM9f66mOnMPWK6AwXRx00qZBZiBqda+oNrzyqrv+ol4phxRqWBdkOabDLJRytkyzztIPaqgf0g
nnRCmnM7x3FflljCTe8VRGUpn16TuQlb29HvsuUNDvOUJVpZYL/ObfObnv87yo8WbDE2kJGP4Als
UahGZ7rkHqApH+7G+Mz21LkD3JV+qWq7sW5k7ALwq6walDEd5KVyDjzA9DZ7A+9aHo9NVIJcqY7O
RYeWXNrY1YAGvzz945dFxCte9+O/7v/TBnYEa6A2s+JOSn2/wGC894E7SEixyPuKm6Is5P4zwqUU
j6PlNV4Nij9jQF/jfHk7aJbkAQpadr2k5LHJtqS1h3URFGXq1Poaj74Dh0AxGttpumxQCZRqYzdk
OeaFq/eNiosavUjLO2ysG9VSgjL6c9RNoFTaJcuhHCZZ5Ss44leP56TpwykAtA4waom6ODYSeJQi
UygknU7V3z1FIND+GRtsJbToDB7cgCr3tp1AJGJD6iQx0LtYxhUL0amkQg2ps+Q20vIiBVgGN3O2
8gcmHvL2Bn3b3DCRABBvQpL/hhfBV1l4SPDpGcWfXF6I2zLlyw8PGFLhiDk+dkUITDRzrlVbfQ4o
DxJA42+QoW4qRB5f+RnjPnJZZHI4JBC4Pn7V7gT4NcXlyrV7Zf7KCbfDDym0DTjQmIwDhuk6Cd3F
mw/lHb9OHgfJctEpLzgQUMI1uVtLrHWUwSof7wnrQq9rZdFChbLLn1BwIsW0ufd6jUCH9ER/sQPZ
kKGsFvP/h9bqAF/St+vPFynXYbV7ja7rgQz6riUYdiRr/SWO+kd6MERsCBlvEJuIucnKpKZzGAly
W3HPdqVDMXyx4otYNoqBNmpJYk370SK9wcCMCrOC1S5OVn3HQFe91J8U/nTRMZupLVYXlIKct4xE
7N1BkOCbbbu5mWOJ3Ad+hpOx9I1Pv/+cSuxwWC9btGJOd+WQqrCZKDGlUmo6fP9s7cx3Ak8tc+lz
CMUIGCpAhm8nEpZJNOA8yibJ4xgBYtpqhBXfMyqvKU3lSSGnzUkBgbLgsSmixNmvx8x7vTN+/G2I
Q6LWYrqP8JpfYxOaHhu1jThMleChg9DNRu/Xlx6t6wO6lDPLBHzDyCQ3c79YxFtrzzE1eFOeBbZe
r9i4eXg29IiM7hUfsI0uPd5k/GIDPuPIRE2YzLG5HX1iPT8CnNHA2umip+iAuL68bWKt001/3/OC
GFK5RFwkjgpb+q+aRqcC3nYGhtiifbZDE8w4fcYwwaO7+IOdx9nHmbJGXLqE0DcGewJQMa0Uovhn
xFcdBGlyfwF4oQt/D9PNPb06sYRTnTd6oQBFvzOqbJfQofF9T6BFX2oJivE9QXXax9JH+R4sLoOQ
9Ans637eOTLMjblXuwh4vcfqz1HBk6v4G/TZExjbv3ZBwgapQ6Td56M7kyFZmhRHgAZvdkatL3vw
vAakk/8Oe8WJdrbWwDh9uqYbxp3S4nwsjhSyjvwu92CJdNIyHoK/1VqyypDkuxwDWFIN7OnjniuL
jJCzBj7Nmu9TyFLNbGQhAULZIzLDZ4jvfNYL4hXT5bWR8WCDKj0PdC7ZyG0KmV0nhh5rS40gH8Av
9shTlS3lttrYso3JiKDOrWdFVfqtmqcJYumCFgXNvUt++kxBYZ34VhGvQCoV1JSMDaB48qle6y81
7hyLBHTvXi6sg8yzI8oxzhxQHxudiSrGhBgi7vmPjyj1wILUtfU2SamFFzwuFK0cpkscsTjWZDlI
Vy1YWWpL5wbXzYKr+/v8tF8C6GCOC1o4IvJHtYX42J4UoUYeqjei4ZaDNZPweoLedu6HgTrXDFJp
Aky7GJiF6Vy3qlu5vJ+p3st8IxHanefgrkSa62+GjjH03RvoVFRq+Y0DQJKjc32ywVkCgo7Ac0Iu
Rdz1H9kT38kJTfVfnxXABOgWptPvUhB0pqpPnu9uE6oz0G/S1XVx+iWOpcHaEyhukJ7r8ObeHdgy
ev2EcYbOdHkjcIyfTgMzSbu9Xz+fsKYLXm046MV5/2UOX9tVzzo+JmTM89e47kErv2liipLlzJS+
amGcsK6CAEdSFMH7H8LqK/neivM7llUUy3WeweEw8lnbeqEDdnpVp7G0oT9RDHRHevLzz6D57F3q
Q+7zmIZYChOhwAAxqvdow/sB5+HIeyovySl9XozDYUbHnt5UPdvt5EepvWw+OfT05nuq5IfbU5uF
kcDsi/AfPV7aicHRtgAPdiXJEcdrds7CceQeYclOycmBcbTkD+0k+tmX3dzf7IBetvZkvO9sCdIt
QjNTV+cBmX7YUM6pYNYR9PXiviXRp6Qmxg2yGYDCa1QKZi+w88HanqyQuubEtM83oTYcdj1KwGH/
9SKV1mio7h/4YqQYvxyHUlXnF5YveLt57rekyLNBH8qs938JK4f2BKl5fuqbX0TrPpQTYPrSBEKN
ZNx5ZmQZDHqxjTrq/PriaBeCTsG+nC6srudwicdZGexa7kg1kE+HpvKqSqMbkMPgKbyOEP06n0nj
bdtCBUlOOEzdibK8kiso8qiGyWHORImJYtKSk4Qj5X1QdsldmxnmE3PpiNRr9s8XlefeSPP1YE/G
G+WYQSRHQ928sEpVYbavI8FP5SC1IAo1TfEx/OVEFRiPH5AumJnOzUpip/lTyvyh97Ces9VObw3V
CQYtt6HqowuhCRbsXN7mjvCDrla4LUccBqIAerzJDG04d+l4rfiXeYT52sm4e2W/RuFSSrI57YS9
/3PzzkKAFSLjIZAvzzX/E4imemrsQDhpFFr2AKbMCnWmVknoYw1Oqp6YMoWhkkHmTWnUY2Yw/4Ow
xA2vcxe2EYCadoWRUeW1c7BgnJL3y5s9vysYTDwxloctB0Y5U9FgCS/Yx+8xh2sCewPP/n/PoYTN
ENqOWe8ILW3eDbgnqF5qNXLgPt+TOy2R88HtVyOcB5yzmQPidU/smrgHEx5iQyw85Q12YZvJ56j5
515j0UYfisD0GsZLw+dhr4ebOCQ3ZreLOM2Ear+FsUAXiYSBt35ULxnFA8+r9dIeBgCEzBCtdesg
MOyLjnQyBuL66CQpFsyJwbRswdlQ1+VMaHwnq/M06erDnuTvB86RFE9dAeyomP8FjVV7OUWGJNFd
I5mlWG27sc4tCaMqIGYrZadOfCcxHYu6cQXuwyFPEuorLXqL+sVoexCGXoBgK1nf+/I4PuUahHwl
wd/j0dwL/55ZEqWWLpjwUfzEskFOVmp1IyOXUR/1ZrRQb7zgln3d1qsghhupxZ5s7GWKyOEkldfN
5WT/4jAPgodHTG8dI3qy3+EGx87xhTiOb7rgTLhiEmBmNBgdurZba485DEzl8GdH+5Y56nOT70BS
/o9O/QPULFN413KV4bdiax6m24ljhO0x9nWclCUw/e8TRfHrOk84AuHKtX8gfKgoZzpVj/5hWkLV
F9k1Psewh4YWMm6JaMiIZLhzDfF76HESz/OT0I74k4esX8d7F44R70VpNmMJG1fBelpSY2LjIkGE
zTu0I/gU50Jt/ljSybywT/eRjZ+DR12gJfIuO4kqkgH0RXWWqcWiml6m33Z/TkIBuoygx6BurL8N
nxnFVgOjAweeNb7XadRdKPSuzaokY+tbNFZ12cRW5HO/mXRrj5Q+L9NmKYi7eNY3OzjQGnRTxCnA
SVoIHSKtBYddRyWlwywbs0lDsjTKrgQnl/JQAzXMtJmBrAub2KKuMX2IvgF5+gVit9I5WOjxs0Wi
0MSuTzZKvhgc4sL3lJ1cOf5nEgXAR3MnGanA5bt1kbk6Rjj3kJb9H/8viNZCMW3/n23SD6Zgl5rf
k1qtJRTGrffXu40NF6PzgDmF2U/6dtRo/Ns9n+2/BcFoaM70G00mGYdApEbgzcRb8hvv5ieR3SvC
BkgFuRl/wPAJ2iZH8Le9VozpJt1XdT3EyeIQLrLT26Jrb9zr/IOATTNbnkhjbKFZqxVp+gLfTvp8
U8MPTyJRVxAUqTcfIYxhOaajmbHzWpAkIsS2XB82n+3nrOalkUahc9b84tc3rc2Iq8BdT7P/OzHv
y2eR5FtmApiiN7HtGHXYbsrAQ0Vbztxa7l1GE1pnwvUsq+YNacz6p4gT6OVioT/8dOo/gfe3+tfO
SCl3Tpf3tV/5PnbfXZ0eIWPmKTHNTVKGA45BT3x4/sEfks9kA3Ax0nATL9dI3Zle9CqiwgYv94/j
CyNw1JR8F0IszX2Tc1WLzfN96fr+wVcYmoa1KjrLFPRhzv/EJUAnPrWJfdOZpbN4PlZ22J1IEpVJ
suKRpnv6XBOUcvEvar9svHH2U2Q8Rfhjqvkk1/x8evJirlScm+hdRDDwOUtaU6SI5dIUt97CL/aX
B5OuiceyBcpcK1v/1au7Y0YPQ68p8sV2Q3eFu8ViyVFTZn371WhvPzkZ02dd8klSb4ZZ4KOzwvnS
zcBbL9sPoW/8slFD2i8SiSoxhq3TWApYaCBwNlKygyN+UZ8r9vGi+lKslb3PJ9QMoWwnaslnbpyD
stwtJvFXJvpzwj3ntVk8QSjkE8WKYyennMiYydRKYh97qUzDL9cJu/CJv7VeWEwbveZNMY8qwBBL
GQvrYCjgNXNoEQgWRCMCZOdjf0GRu6MwR0kaFN6shJAajXt72LMtWiqRt47P74VvahBR3fXvnwY7
UlbExrdi5sdXSNkCD7PEJZjESogyiPkMH3X7skQWKu3LlOahhqaSKMH/+X6pYfn4g2vkBPOMFksb
R4eqFINja3ganFyKCrx37jp4RkQ6LHhFBJZaoWRggQxW+YgDUQ9WDbReG0nVb0pQJpsXjfulkNTZ
nXyW63J4Ii1m7uFtxtwTGApDNsWt3bfNcJRIY3b3ulxnLd88dwaQODWaQOk6dZTMF/FGvUg0wJy5
G2AtOS4t/5KnMZgfwxey9n0SwKHm3EdQ4lJFddCAKfQnxmp4a9qx422Y0oYT4UInMimcYl1gyZ41
tY1kSHI/q/GojsnqGr+4nkiA/2b6fSSUY651f64HD+GdxiXUP/bJnUFTv/1wiyxFRYsASuF59wcD
1k5ntO3mEOH38ubZMUmcZyHliHxy+gvoxQ7PNt80NuquW+Wx/Jm54GZwGP//XBdCBqhOT6zeRLz6
vTGWu2bfz/gDouB1K387Cq8NmrmL87prxLSm2chcap5McC7dR49U+MRgNKYLogIZ/4GgGPx6aKfJ
FIsj89gAkdfQia81/zCjQ3uBUPgrDwUQvnJSOvjT43OUsSrt0kEMx1ZxM2TzbgFqDIWti46KUpr2
Bf5JduCEQnfqbXPgoWZaX5zFOQCCjFVzm3rfJyv6rLyiFTmvlff+XhLkLzqvpYe+UJ6/pVDr/9MG
NplGA73vPv2uUWxbtP7njFDeRIt7+oV3lj45pf2uy3M3VBcOg/aGPyQZKlH8b+IG4G7QNk99ygV5
Fbsqu+kTHQxXMzqHbUt9W9wHm2N1+Bbeww1aZDZztULRQuTHWuotgQYqPm5Y46BiwhnPLX+SsXYh
s4pyLSiPXXlL4/gbc/fOi7F4RlKRQisC23yTBq4JOJrGm7HMQcMwK8HNdavWeVLCdb3RtoB8YV0o
urT4k52c2a48WNwIyY47U2qPqPUUPLy3bpEoS5gG/amt3uXs1JFnuPjGJLkeezM69hT9+TFOJnd0
2vBQ6Eg/UenQ6G8j2xogsQIxeUvvTeGWgfQGlCGvDfYhPR/xchas1DzEyK5aBdAPeJP5iwnhqbnH
A+CHWN/DlCY8OOTXLUzy9UftaiwE7QJnB4ghOEw1gZtr4CHK+hlXhGSB2d/m44CPjJYoQRkszCIu
+0LBVRf6XX1HJZ8CadGMaOb+7/z8JlC0DqgzBs0rXwuiFB1n1voFZ121J+AQQSkZS0nNzPS3w0EQ
GzZsyS7qncn2IeRhzLBgmtPBa4z6BkJw78RjKqQQTJLrB9BKDimddJM2bP4lvFDxh0cJxQi0GT/Q
urbsSRAxqLt7cvvWsAfOTW5IeTBlqmCAv0lBvviMUhaoQWWMIUdaJJozH5yG/rJaVoQKyPRiOl3U
KArnFmy/Nr4/cQo6ow7iWrsCGK0WRG2FI1pOE0C8mEY7wBaF9DqbjPuAR9xHvGWO0S997rk7O+TX
1o3UptiQnuPkslgjjDfnnYrlvH0jNlbgBTrfkqIJxD2dswzBObxWEpU4rbncwmbrwyEzzVW81Y3K
kgTqUDDgyekFKFUOTT3He1g7LNr1dkUF3WliRCQ3W27R2YAsfTvubK1RVpawp1tX2UkmapY9+Tn0
bX4xalGDR4jBapt0flDworv6/V4ym42GzNK0BZU9gxsOA0kWjNr8iJqrIyONzZ7bwy8c8kIYv12I
yCEGwOK5iO8jZi9kpfvqcVBNCMj+Nv/fc/KD9IzVDF6zu6qGwE7b7O714t9hCbXX5irbc6QyqR05
1Aq7A6xWxknKe824zp+trgVHcC5fmvj2IpAHJMEDUVSzkZP7T+izkezg7qZhNNHbCAf3nuODCaJL
2CO5jtiXiZEbSlbDMmm9fWKakLnNkXr+72TQRx/I6YZJlr1JrvSIDzpWVVuTxkrE1dFkCdzBuhad
KEY2Sv4AhVIaAcmIapj77ICalQ7OxcmECYPStYvfMbrEYnMEAFW1Of/WUvtOyHpIYINVcvr5nJHC
DZm7iL5s2cU76cYk9UavpyAstUS6mGdAaE8ZTal6udeDd4wGqWxhcNBrTpmv1C6JlmwfE2ujD7wA
lbQuy/oTYvvNqQfOvUnqdjrw161ddWVaBgeF1SFhiFmGVnzOUg0/PVQ6isu8pUZFFCLzruj6Qv+g
VeuTkTcaynt1OacTz3Q/RjEwdWqJ5EKOLQTTGVNhfO7zCWyEwo7/ZYAQIN2iZnHEbwcsftSddh7p
dTXER9HwxExLW9WUJeGZJgn8e+LiyqHYcBJEEyza8+VKeDi4DufGkuGi+dmdJcx8abm00WZIiNLs
xm3m0BGJH9uTdtsHfVgkFVyZvaynbkoxSiRFOT/s61mFTA0uqSsmVQ3QihpkB/BdR5msa5C5yJEG
Rt51u4Cnfn1mFWD1V2NsIf/JQSy68/vmxkwQq8zYJu/+N930XJEczG0vEh4SnPZ4KoXGH7CO1RvR
Eksy1CgxRMX1dLleARu7XYKzaBz6b+z4f/ycfYecthhJSWm+nBW+iMmefPumD14Np3xtpFOgvFKx
YBO2dPALSWltPLV9BzpafTNWDCu2IrjlqJBrv7XA0Di3qkWSpXR8rCaQi5fVqbZ/AmDSM7L+lKzx
PJS1Le8P0KrzeNnnU2iZHjdBkKuYahcxtmlPIu6Aj1T87Hkug/7hvMYMtB33hsFP6u56VVsaYqNQ
1h8IQ2awT8oC2VojfGPXmd7SNuYl7NgAAZEyAievdHLVDT7mqeOJyUEGadeeqgeYbKZdBx827pIN
btXXshfEELHK8V/RKFT6/7bJv9eqQwOE4Aay/sWFCdH72cDvuRMj3rFMoS7HgPdIRbMOWjoIKBhS
F3ISQOPADrWuwv6iI0GDPUHIYRIe28AjOwk17xj7aaipUVeleZH/Pn+conl9d7YIkdc3SNiUuIVx
4ApqOLtqR92cB6QnxMT4tMWTNYcCJpXUeV/IpvbpSVEoLjzZx85RAL6iZ7T0OB5zjFpoMZp7EXDG
nl1m0SGJmnah8/b+ws6FHFqO0ZxQ/ito/t0QulA3bgDRR089MMLneT04WNn5WWaG0Irj/3YXjY0v
2M3KSA39ykaxZX518bK7IKvRHCP0Ugwkh4YTxfLEzFzSbu2GxcdEd5jHqLcdUHxv4mpNRke/Vv8n
AeolxqZxIMOc9qVXRM6VW/FGmO13cVEUIkUd7n590lAXDSls9tXZ3OODQkP34MmfYC5p0g6TZ0H3
Ucpzh2V9dpX5FX3bRoO8JwS6qcfGiwRP8+AwPLuUMux5tMmKbUxrIervPzzfuiiIrHTpQ1Ro1JSJ
wHU5PlvtzRb4EziAsoMhlzsA1syB0P4erhmtfJyo0mxz8gWyauNFYw4/x1kkFmD0MCcxXJQORXYk
Hnf8PTIQKfS/tjhJSs7QKZ0Pzl6dmLiDhViz1/y+9Zym379vW/vZlAzR7Cg50TWUptnesOwvXKLm
+FPwZNZ87CRRITHEbDh/cscZMl4W4ULG3q+JgcaWre36y28jxg6EnFpO/OWUoSxEX/lq9tIL04kg
hzTs/NTrnhjHV6MTES416n5Zy7lFxn66hIGQTsMvSTN0yD1Ixtfh9r3R8jB/uPWrzy1mRYl3Eexf
phfBhgDEr2yCFNDrZbSDEt8mAZZhu5SBbmaYlcom+VQUv0tz9uH/09bH99ZyQHtvHi8HQ8sN7QC3
278/x6WpS1PibtLz8pIOi9S4E+GVU7s0Lbj9ZsIhfFVSc67FK+oUGqRomFeIpbnEckfs4JAWpZ5Z
F0ekOKkSABvyR30RBAUNipiOgiI/yFtr9RMNruuMTlDc23WK4SLWef72M5fzskWYigyMgBJrrJJA
p+9+ukykY78MsPX54Yo6WElagdPDl1uWTurhKMv8z9g2dI9vp3K4IQ34yoX0MKsZJ7TRgQp1QUvV
ScpS0K1ufXhSj9fNwP+gfvEvfCc0BCXtJI6h4WGlQK+2KHsPPa2qtqMydhsmMZAl66pA3mWgJ6Bd
Hq27iF2R1v15tLvmWybCXLMMDL+qsXg7ScVJFobjcENfKUAjOO7kTjNd535FCY5JW2uNJF7uJV5P
k7zfC/66czxXNgZ7LG9wntYLpml6gLoYZtLOuxvFcL51y/ia46/yWTfjNNG7x0FO++3rVi/RNjf9
m5UuCpPMKmDb1nhQroe1hG0+ffcldu8nLfQ9qaG4vgGcMNsvnhl2j8StNluJGW0tI7j5kPZGXCni
hDx325JAlFolrosKGk7kq+H1Mv2SrI/nn5Lsirg2IVk+yTLwpwBI2AYpi8QE83Me3Ps2VIqbyHzy
Pmbl/QWaFqKNS9we1SdEoR+5R0HQgp9mrDDx8savDvE8wyW9SE9WDdyrZh7pOoS3g9CZ2tReUCu1
ONoRhbknG3XwkAxc3BboPBE3gXIh3dP74IAX5ceu9wYelTlIpjFQaX8WotXGWh2uVABTBwZd13eO
IMi+1wS2OdixMnFn5dcmP5DzQJG72Km9zUjhQHO4SyiD5bgSzsoYvNrEq3OPs1T92II/WDmfcluf
5A/KRz77SDfiMFYg2YUHAQAafgC06Bz+orp7HsVQ2ECvCyQBPXz2vb3BPHjIw73/LMgDwODnVnts
TwJr0w9LPfq75bDMjB7akRW8hyZ7g7qh1/Wf3kKy/0LFEQWFJ4CdZaGd4zvym1oSdMgLtdEmxcg0
RlnZT5zkTBcnqWCyruVKbvvni7hRCWS4g4RtGeUimmlOifsY8YS6qseBt2WKL1lGmbsuyIXL2cfh
P7dvLMurw+H+o011xjTB0AIIp55eHtC+XL58xA2JVxxPmR7ZD8pP9NP92JYWb+XJQ0QZ2RwXG4+Y
E8c7rLBKCS7oDA6CsUr1tWrssd8wo4Oxj5QSlUrSQHiafqAA7+jIAJh8M1XZLTnYG/OiU9VBxwMr
XPZEUkNWRPBddQQUKrGQrUFTSLyjBcyejm2/88xoe1zpMrXkh16XJmlmoot3bmfzJzpXkxC+9pZ2
OwztJOrh21aPqJXkScpOmoRcnaHflY+qRfDLr90htMEEcDBShjWJbuFgN5ZuE4ezN/EgpIqeG1c6
Y7yC4sqUV0r3CA7BYSGWZSLybJN9zyHduEWwCw+6MNXPWJtN3eh2CxbOeO6i30yd84ISfH0thv5b
wy9PpWvNQk3h3feXy0imkVW0j7ypC1KXopRG8RZhmuXKpbDetIitlSgdXoRfhwePr+PcX5RuQkPe
6lbXzfDAZIqo45QqQFhKCFwNRzajkUwUK3HHG1MQMSQvJdt8c1mISRDKcNimCpWTv7mdFX3hY9XO
bZ6oBfVn7+uGioJHtnY7rc3bIw4vOGEpo9jNKvWzGeOYk8ITt5EVkOgEhpH0YfWhuaamf4w3U2QL
L08Gym0u+d2kMuBt959EJe/B6cKCkzuHpAMLWJol1rSXfTB5xxS20p3i+WR03INfLZch7IjBLL+h
P/X2eJ71aruUnNzxfNDcd7J05WgrAvZJ2kblAIBDsVk3Yq8tNxj2OJ82gSh3OvdJ9nHfFJKunBdE
56nyrhLIJNcNgLoGadFaNOghBbwOj2WibXLifKH5eosS5ukX+AOp9x24u0inb8haveZeeay6aQ26
DNiw0kP+1nfFoQtfB2oFLF1V8k4Y+KDNl3WnXh/XYa72pTXkqY4dwgU0ysE43BDHuRe+NTITQXm/
IxMsMHWEwdLeGNIAIoH479wSeAx03JBaoNgAvkyUnaDU84nlH3OpPOIa6XM5EM5KudS7pOhch04R
G/kJcnTPFVqfXWYw944xe3V+dpGRtCIBjIFVRpqiJZPdPXGta8CKxzoETDCPGcIJDQZQ6uw/8yow
GaehxSjhJ/9id9nFHc9MRSZ+c1qIAoFE8fSc1WFwqkXWgbmSEuGfZ+baFrBXnHDfESsidBA1C6ZU
7DPqt5edHnhIArhlZ07/upbzyJVIILxIa/qd47/JE6vhQOZz8es9f75Zb+hBBruVRgFcVS6gnyN0
+3i7MY68IrxByTD3+iWYX3gyv89jrJ87tkrZ9Fqct7e9nj/QIoUAqfkiHYEuKUQBzYcqdN7oER+6
9zcQrGQ5QBWEOSQobSYLyJITjDTzSgh1gzkDFV/1iS8/TckZoNSthDAC85fyFaXPLaDIsm+BCaE7
RgH9cFHISFu6C0z9dNjy6yLiHEmm7ZiTTDl+qsdaNp02P+2pKAnCpQY7igOTLtIgZhrSfCWVtEHM
Da0CPxDLjlxrWj5aqlt0lEdWIlrKqsa6vZIN2kYqN4lApFCq+Cnz/mrcRhjcp+M/msZA3SDPyCTN
tPPWuoqGAlWpdArYE/p58YKdJ8hWPVa0XmCwmqKEdyV4EJChHBYpLjzE5BcCxRoDVARuKniZz0h0
NK3gLoFjjU1J8HENRlJTWWdYMDhf2IIjdxu3LhLgkbFnaTpVJDYLZwEIlDPQx/Vhgiw2OY52NuSf
dBdXNlEldxwQP5P4HQ3S63DnrJuZJoMjJxhbYtyWFZe6Xr4P98tBrujYODD9ZHcuuOocDCrWejge
q6Et1wtsHFs7yQpQboH4xYM2CaZ7JdOR5694gemEYtQyiZusc3cejAeKr8wTolfYcuNknEl0WIB6
caSBjhWIDkzzf0Wa9F1exNSP/nunR0Z/Fi2dcuBuUo1tAJKE+vxMW56oY4dAkdR1M4C7psJIVTTz
pXpR6DlPLNNs9goYZUK0IiRlmzXUTLAOYcvXBQQplelZaIMNbEs6684AJjnfZrLOh56u3CKfgGK4
nzRMrgW94hBYsJ8oCgS65FeRFXZvuhF0lrdGRzbRaUGRip0N3YAHnCQdqUCJg5iK5p7wbK7rHthh
W8errO4gN81qiSx3TAGLT3NGMl5dhhQsG1MK0sJovKbalRYoWPXV8rQjsL4ypDQOMVJFxFVczEIN
pa6/YNy9G7zHsN0F+VesQ0SDh+MwdGFN8smVUBI4Ls3eENduo7UoOORJzvaeLZbFBlJzZzhqP0tO
Gm1DeWp1rT0YrQZx+t1IlQH/XXxaaa4vNXheI47hhNWR4RhfgpHt8w2/FuaMSHLelcMd+crStp1+
ulx+EXv48XRP4tEpE+Oq+lJbUVD5+ff2S33SpVAocBK41cSh3acm0qbTBeRAwhs6yL5aYaCyzajc
oob7q132+moRkrmsYsj1nyJqQz5JxRb8AVJ1wqZ5X2U7mNflxqIaEB2izDj/GaGApLrBTmvg0Z7S
364Tf0U4KR9bNmU/L1jPRQ1ng1TNeug0TmfUg9zAzqec11CuF4KxtU9f8dNS0d4M3JqJv+FzkOq9
yILksObSCuXlb/sSgAGHg8GeFAmzyzmu4eorlRMLiFes9ZaoB4lUFFp/uE0hKk2JjAPHytq1B974
Ea2CyR5FSCIZ0jurEEoptBVGVFa2Uuc0L9ib+BiSrwQruazlKx0kFqzRnHiPAe9XH110u8Z7pLLR
q9ARAbdBCavNBV3ViDtsvQnN7N6zVN6NBe9B/JCmNWpK1RdAvsf5m8WxjoSSrIPBFIjKR+48FmcW
TOgQR/cLI8hxIlyOaVJG/twd+dinibz0PbIlw0QrU+JlnrOI9xU3dUe4QviQHfy0voM//gqtHPMI
05zp6u7MxWl865VSAZlGnOt3gDKn09Q/U+GRUN/2cmqor2Qg6U1r9Zkmxu+FMeDq1AkNR9X2jGZJ
Rc9hB3YAXfRQHYclMa7oZWnwr2PfkBspTeVldQNp2LL4gdqbYHOffDQWZyUyUpguvl/UJtHjiAiD
OfINzYn/jT9M0zX2Fx+uMybA6utxkTveePG+PDP3TIvpL1PEl5MN0UIDEe7hyYayi7BlNuc+PqEN
Lfw8qFEq4+tZlUbtq1QEPg+yHxBy+B4Nn2VX2z6dOL13/iHdqb7bbXGknXgCnIyGXzjCcr418KcY
ZN+AWxkX2+Lz6DGyGt+34ZU5iNLirGWeiBttADxsL59S9PWTTtIaQD8i1Lic1r91gXC0hDMrE/D4
UdNplWIMBR/HEUtPdUJUC2xFxIdHsE/BJAIRgMfkhFNAj3PrZrCWPsvXsGRIJEGgJ/uXvXt12j5I
ekCLi6YeHQnpxhTx4iqy97gF0JI4Kl2OWVyeCPm2hnzuV1vf0yrcAl9Li3hNpy7Y5EzzZcXw7EVb
wLsnZgEGn+AWNG+QNfd3rodQCaGJvBZlIircsL0DA4a5bEcYoz0e/5ony+RkNOU0H41rNZCiSw47
HNcbNQ5KvZsS+DiMsAktwp4w6RvE0yr0qJIDU6eGOl9we/gKIIrVkF8RseE7I/W5EMQjCRNOO0EE
1Z2qQe/Ge4rv5D9VxaObWuhMUnoA+ST8LAXkNeMfk0DUszXBoIG9XbAJ+wFtt7ysCobQ3ImMsmU2
f5LRWqY7Mq4kOIu+o6TWB69+wpDRkxWGVAj1LpiOvY0zgltfvr5rneMU8FuC0dIYVAueqsMd5vld
9c3W91Pk4oej1G9HbPWY7mYrDTbucJh+ilv6RUFbwxbSwLXn1O6o/St2n3d9loHHRWFWt1wp5h4W
SosUNSfhS0Y6EwcoaBov4RWO7TLuSaiQJfUfBZt427deH9wEs+6ks29uaNdy9HIRxrBb6xLQCkN8
HufbWnenQf3m2u/5y5CG+tN7zxOHaprdMBCC39UbQQ1RBJAQempvNykFxC5lbJM39hWzLYcLEj8l
bsei8FeRqptcX7JspLtdMOUPMR3mYh/zRI9qGwljJHK5UKk3Lz6qi7dVHYDysaDJVnd4UPYQBylI
0Sdf4YQtZeLAHi9U7UoSERVSiHp185ZuNvdSbBGFM5Hyi2BPXNpR5aHk5vf61vPJ3l4y08aRAEbt
BdBalvCO0LcwOIhy0UlJAJHDfLnNEmJ17P7XaqskcfQ4DOTge77TX5zPLbikkfRsXqImlYkK6brE
zqfFuVsqz38qwNrTI0P7QF7pbfxw6R1SqbG55Vwbx727P1K0+ygJka0/YqFSjxd1TXFvgJ+M/HrP
GqqYh8Z+1Cv5/+xJHTs3tFosGDbPVK/FrDhF7SOfVgdwmXWmjrGaZyE3m09dxOVKLxGgLOQJDTWx
TojOfSD+9K8sye7Hg7MwKT5Ac9G+98ypMY6jGfljxTL+U15KgTELG4X5GV1/x5rj8xhY1QRgwS3U
jo4ia8mMWuenulLpWTrrdZYPikv9TEXH6vc86WfPLRemXBmTYJ0uvEivkFCotlR/ti0GweZ183t4
GAkDukSlrcB6THW3B2La2tlnmjwslmqLZIYL9LwJltoxMLI/72xbT8eCk1NzYTJthEHikAqeeuZW
2lVntT9gxhT1BohPh30KHCh4u0GW30uD/3T7ZmYn3B86qDib6mBmhXCplykWGjhxhT9fGpfIjQSx
6ngHAZq9QPVCZqYYGRwrHHefrxcejXPV77+JAZYJNjfKQNoslccv8oFWA0nlrNWUi4MzJfy9Vjih
13N9VntJu6qDPeWYU/CraQIDijJ/nnKPCB89/vfLt1SU+aIKMi52USOoYVQhGMDdef5o3dv9LZMf
5pIL3A7I1pDenXWrSMHBDYuK9i7Tr32SPIYy/VRAPq/qezo12ylkGesqf+rgDklzAQDm6/T5qvaQ
GcecGvVVdET/v34FMfyHpdcrJ4iB1PwAOrz0U+qLAhvf0Pi7ElXNmOTWKBgxVM/vW5JHFI1efiTq
yOVSkh/cJ/YetnUiwlpvYxDcTjFqA82L1RqbF8WpD4V/sWd0wSrYwnT3sZJg0VaQNtorUAZPpc6+
9kyazIN4e0T0j61m8HExKphQeK3yn+Ce1iYbuIIMd18rXKkhSTq838PH/5fXu+fp7nat5RKYcXGh
XaYL4r01yej2aPlF/jJUjXg2i9bdEuDTFufJPMM7qYt382L4ZK83eIEFQ+L84LDcyOKoRzivb7vR
9fdUm+qE7LwYSSRXpb+0U1MnQ/yOzm6d1DRk1we1k9wshuMK04I+k+nW78EpmiYT1G4ccdgP9SPq
EX3S0GWTQ03SPhhkUWsdiqTjHXZ8Wqm2gKuZ4Bz293NnNSr2sCABRcjj8XxM7Yd5MMmynrIfM1Yr
s3e3sT0S4F2c6PNZF/ANZO2Yh9O1S4fsxrqli8lfIKl6wlO2gf4mO+Q5qcES2MEkBOD/3PVot6/Y
MZUqKPuio779qjUJU4TPu9g7h8hcr4naZzd8RN1ZveV5sXxrIOp4+HAU9B2Oc7cn4hCIqb+yNJGE
aHKaAJWHYnBdBB6J44kqxdxPDScoTNUfTaHtxCtmh2dFg/5n6HIm2bjhEGVI/WLovP1lrb4zw2Zm
uZHjbXfQKQh2UVGTN2+LvYeh2gJxtvKPWF1j1EZctq2OUK1wXDp4qRG4L8sGAE7bgcWjnnlGyfY5
gvVmYAudJytXMRRlcZQ+fV8DOU982Yy39eqjYpDSiDaQTqUlqPg7+Iu80rrr22ong6zlSlexxH0p
EwVArlR+C2pIedylKz2+SErYfFc9Eqg9x33m1VRQcNmp1+kVRpyjUG4SSlaMQgXFd538z9tZAOck
rROAgAnbrHgHPm5LMcen9AFHojMHYoD+MOB2/61tTpWey0u0MUW+RSFg0IQ70IBHhLc1haDz6gg9
auyiwOnNmSv8h04GKZvLdA0IA60kDHK9EwWXKIZDZx2JX6FZBhTb/FZxMxdH8NypZRh8r/hMj9Z+
WiyOKhUiJYQ64xj+MpGzFa4GNGhXU2i69m0wWPUQYRdXuVTcB0DiUsWhzyli65hym0sfGR1yVVYR
BzXWRO72ONUhVM7b4seIPEtgznvDdUYrh5c0ao9txoCZfDSSqJZcUdbvSRUWC3l0itwAVT/5mNnJ
R/AkxNMR31EM8IcDu1wdx9ouPUJJk681nyehMek3X/qhTM6DhfkZ90mBd1hE3YQYDTUAzhSv0+K4
p8as6twnE/994ZIUYhnOn72YKWyAOi7YR8eEqWWbtuCLzq0AK/hWexu4/xGcCOUxN8BFo3woWSiw
qNqePCBCAjAocuTunyXodpKNqV4tQ0mwWX0MUEChmwL9LZsklkONuebVGB2yXbDhuhm+G7af8mom
WKZTV1c0TxLpvDUSomBoAGAffZEFS9ol2hPN7NnhUgjPBxpGuX0J0hXg0KBGScUK3wmixHjtVJJj
lLjAFBSoJV+AQxPPVma4lfz6FI0bXD97mmjZE3OVNu4G0vJ5yHTGCvN3OJrLDRMBmClqug2SpwUG
tFcUFkGswRyLXM5bhmb7DDvgShhrFWqCWbIuWs8zFP/sCyZbR4cs2Cst7W+YkUeZIFcg1RMafjgz
QNtVnIJHb7mIcK84xpQwU2W9I0HN8ZxbrvJX257e2ABPqPQdz5yWHIHRacrWIYJJ90Pgd/NyOWp/
/n0Gl/J4OXeWz5+z/zKdks77A89peWLtTxa4jzL7au3k2jTrZpjYFl7cbhIqPWb90HGB3254UB6z
e/3YjzLr0TAVstCGx4ykLn64uSAQiHlC8EGJ5SXCS2chOh18IW2H0RvdTxXLqyPTS7H9/sW8lPi8
BNua3RUxRCEJteVcWRaEcUcpL/l66NOU3bpcswuN1KjG+OCdZLAviXzCPjtQlz6mXnxgYS5J/sh2
TpmU/yDKL5EOsizR1zTz2Q+Um/ewEGz+SNNXIQPtM4IauqOG6iFaOWqx7o2JIyX4UEEKXTYJWB/w
dJLeb23QicLyZX4iC7z21FrgrxKAKjg5qGd91hi1/b74nGivq8JLaUtNpLQC65M+eRSmP01k5LVK
JNhPpn/2TAP/cv3TC4yyN3jBFIQ/hxXPy60ktP96qJhvrfseieRJCo4++2n0+fE/3ykHnW8bbGdS
bKuPQVWVS3UEt3BeL5Q1Iv2WRmDqI9hUPGpFHT1RVLRzZiLvge154G7QoQFOesMBzUl7FzzCsCmb
JJiEYr2a1q8AEKk3ltv+1uATpYgF1AG0u/J3Lywfly3NnHZm5qd3NM/jZFIVWU1s6Gr1DPqVq+OV
28QycXJpfD5tSIaDpCtb2F5r3JLxo3dxa2zZaXsSmwvnyzCm6j82b5rVIMhxtSIemZToxzfyBS+4
nPynCh7uV7qh9a595aUUF7ZQBjBV0MyavaN8Q/8ygDwRSHPShQ8xEPfVUYa2JPVgnDK9vjpS0beA
S20zqpFZv9EI/uzl2NIm/NvrK4i275PdeHKV7XGLmHo/N9Scb9Rm3X+3FJorYC8+zeXyxcpr/req
ATGjX0O+TT7GElbaaretYD7D6MuCpU5NrMbBbgxyV9klG6ocSyRvDSMbw3KfJl9fuucqFqWE+zC7
NEuXD/XjSWSx4noeFExQLuEkXjLlTAqMf0hhb7Az/yeF6H23uOPjg4NIIBOJUc5YyZunpcjtjv6J
htIw3KyHsdiG4uVQXC1LwocVVX5YlFGflTbERm7WLokHnXtj5AOR1+IO4udo3HUEqWr4qOYTaLs5
3UcNdu91ls9xsl4LC4LLaEoqLFvPp7HDIg0VSA3wVmGg54tiVmr/DGAhsmrWcruyp25BPxlnFOKY
9wxZaYHVEnu7rpMHsEzrqyHbT7PTDaCg32eN2lXLi5ZFy3TPevDEEQVziSQFgWZ7/lLCZJWAIjTf
NN5eL5184g1l9gBRQ2BH2kNrLoqcgfu1afBfLK7VTT8A5ECnKu2XKA0djRFW3MfukqfDXS4JXaTk
A8tuAhxTYD6LLyVyPTfs7/4SCcPe/JkLKUFca5TJZs6Eg10z/1dGEGuqIaocJXmvgrGbjP1bo4qa
wt/xaDtcG1JcEWIscwXX4fHqKT7bLaiV6Bgf+2lfLF0iFhcQFX1eHEKShEedXEn1GcZEegKU3uhl
YeMKjwBdpFX0WcSCY+jWGTu6nxByaxxKZvHi8my+qzLUITCefR2h1LhW4SIsqMd4q4PK/AVTcCeN
cBDzu74ExAoB6mFKyjeBQfr3Kv8jIlrKV0aFBW2iLSx3k3Nr7ZvDWvHyZJedJIdwSEAUY8wuwkRQ
jAV1lZnidyEs+GBEfVieyeNM9B6200902oEP+2x3aXIEZCgVLBKQXxP6a/u4/w6lkmGvUheZVWaX
F9PUmysKN1UluhE9HhRyXgGpFrRoNpMPUH7UIPpBLlxZvxvMD9GAXtRi2ar4G/wNNPTYM7WQE1j3
+jOwSkYqtbICZp6xuAuJlAxxGtnSSzf6ykMOm7L8LQi8l3j1LYam2BCHSweaZQ7sTqlkT/s6Dr4E
ijQ6LS1HDIger/bniPooW5xPy2Th/R1NNNgQir9cQmjcIIj30mahxS6XG/FagxRV5NN89N7jqqhc
Xjs1MoUSI07vwwGYbNpo6C2jBZcBR5JGH403FmDgf2tUNdtpZ1G8EtrF9OewvaFLc4dwAoB8E3Kp
k8Yb94vK49NeY7ceEUhPmrI+GuS+Me7J7TH1nxp3NtWTogISKeTh//3OWD64ksWhk5NBIDzTg9KF
I+QhI9q8A3J5/+fAQ5ArC2HDnQPD4wbVc1tcQQI+DPnatf2C74mHERsjHwk6qn7jenLvXs+6xj7v
AT80Cz2zTUY77g/pSJ3nfRLtoyZNncfGOR3i+RFtKerbOUO4uiOXN8w5xilr9LM2Uk+QDb6i+xjd
VmJRvZ1CizQILQZ3nVSwFy+r0t/gj1Kl7OXGzQCA2cM8JMwBQZWG2T6KbHPCKnjuAkdEzwUP0wJa
AA3oxvtpP5RJGW6AD0mbYIa9cjYL/04E3Ii0UroYfDqKeTJsZ1jE7DtscCvYUAg3QZcXcOgh7Yeu
zM5szT+KNGmX8QBe+8tojGHxnPtS8xlEdsYHZXfqfEiD4MHlwSswMiGcMzmUiPEnR8GvUNXudwAx
u1EygKR3P3rkwsf+zADkpaQql/Yd+0SuGlL9CV5OGEVv1l4z3cNzfsxzvnErIyHU/84NQBPsZ8KD
KM1vf5Rt5iW57X4tbxaj7VMI3Vmk3bEeIqym3+bDisHqLOGnk3h/wBbaJCIhBSFZfuTpm4mFz74r
VPEowb589JUraDd5JJo6Un5YHRalX/RAq7BQpkNZoGVf/+BUnwb0yLhZn3GJQGFcQpbM+vd9j+lU
W6G0EEnqDSg3n6XbOvUQuFwShRXnvup/Z8b5YRMctc6wmli9UrlkhKgofNLD7r7d0xpmPEDWF0Vq
Bf7pHoPCZfV1bQEeRmRaa0X/yt5wZIEq6pr5zaZWY1c89pu2SOAtcZJ/YUWaJWV5jEzjCoWJhS2h
yava7d84AtrJG2+QxDhdkhsxj8ntAaPxUO6oS2KWGPLTwZIpDDeLVU7kIeDGsWopFeV+Voz1aape
rCJ/Fv0jWwMLu+40m5BdRUkIAauEl6CP/kFdlHWbFdnby0mj8CYKJj6iKj8yFoVmTJwvY5O2tcv0
avUej4LVjK9N+A/eHuUI9RReVXUP71CvLzVS1qwcf1mb4xSD+tDSyc1MNXTUpG09ltLY3zQHh9yx
S2nZtdt6fVvQzN3beYfu12/jXglurBI/1hH14ARXw3r5iK+C13/BWl3fNnRzX+zyX1IE4AQ30v/m
dY7iO9lF1dbsR1lyPHVUHbraPNz28EBvalDH5+0zbPWoUmqEJvytlunrhJMe83CvsK+vVmz63NIP
WX/M9dzdMmUjCDqw+vPku66Wtasnxn4BGiTmELEGNEriMIeahA0zr1EH74BS2vyqb7RYqP/bPMT1
mr0YcyFLa1PEsEvaeAStQxHRrMXg5jxXyTbVyFBJUas6S5mam8vHWhPK8PN5y0x2lAe7PT/kQXiR
WSeIqjI9KgQCLQVpTSB4EPMQV8yUolfBRSoo/s6+sTdW88ngW3VEf0MO9I2AQuyx1fNCYNeLj0Sf
SPGZ1WQMa7yd71+FR1pCHQju6/AY9vIOpg5zN/96gTBb8+/l9EGKINf9VIN17vVl9f6ecSGmS/eJ
gjZd5UQhy8UwD/alMY6EURkoSBENp0d6HgXnDPOYI4M6LC/maDHYSb5V/AwzkqUMzEJVQn5G9mp8
eafeu5ldZipiGcsLMrnz40j0RbSbsvFkfuacYavLe3ac1mRh+tx34KqISQx/7KbEYkuTZcAw0lft
5joTsTrj7cU6/877iJYj8o3DyheqnjD6/JnpEvpyaNkEytQ2RXJ9O3x5JoIA9JRHAhLtyAxbmymj
/wrrXFma7tuNK0YhQ+Bayb8hPD0bIpk3Zb0SkzIAukWOCCsaDJvrZHVyTj2xbRTn9UqV/Dyn7ekP
/HdHXcMY89kp1umVjR/+pP9S7XcnfE1JVwn9xz310trkCwBEnljL82DF+R/hqYW7wRFtH9L/8t6D
fBclAyCsIU28X6gozfmJvY6QeoDDgmhu52aCWo6sUuJ6sLliyBsFH8U+N/OcPrNDIPpu/LTcnqwV
gpGNyJepHMAkT1WC33wq2EI+fNfQUpt/4Y8298eG22TCvOSJYozBT+6SqKDSmZootLw9XKDvDUvT
dwXvc5B8fvMHKu7o7IjYMr4yM/SFacKLb/1GqgEGbGOIEIwbegSPuQGw1mNymNK38gH2EPtH9cHi
QeqsiDXO8t+S8mGwWkD0IcNlutVgtxdWML1Z2qPePvrgP1GxWMR5t8n/8tbxa8DVLLYTp4eDtcsg
p8LUAwJrysDMYPfm5xzFtYNmm+fiWlF4WYfw76UeFGLZDyxobDc0X87tKyS4yCL3vae7/d73sLxp
XCU6ycgsdL6SNwHEsVJvGMb2Jl1SqxTqYcCHoEXnHHyQ6/GoUu6S8o8Rm5YrnktJHE/I1JJbtkBJ
rR1W+QoJCRqCMz0C1fnWsazg5nLbxKYz8cj+IfwB5BznHQCe74BJ2olo7anu5RdJf9d4wJfs8nQp
+A7ptLuNutNJjMuWeb1uU7Q7cDwf6Xe065uDLEmjm3e7K7I4djg4Bb8fJ6jO+kQu0Lz8uZpe1JIO
bSV3XNVAB4d/OeGa4B62uEYLJHlg88DzYPM7yWqGNjLvxhpF236QEXu9rlzwgY/6q3snykD4rBqZ
ViQD4zLgIAGbhiqZ26OGg0GO5sQBP7PeaX5pGOnVGsj8XL+Yo28g3lZ84FSsDyCln9o8CptNkINJ
czdYl8bP6fBGXpEt/aY7j/l/R6qZbN2PLAs2f9WB9vU67FgRlYR1N0sidXaWVOvE6f6xL33Ht2ze
0i8D3LQZUc4ijrfb3mD151Upw1zEjIIQeWcmDXrou2eegmXqLkxeTW+SKU+SXnj2tMLAtOripKx0
5AW9rkxFNGEkqNLVYYRBF67PtoT32Y4e1y5a2iu7GTFIM+COpPbkSxiAMK7f33bjE9cC+KL0LGPa
vWt3VDpBnno9XyLIjBO1+9x73BXMTnirMJJL9g7eFDXAJVFCr0ui5BoCb8E9dKTa8EgKibc4DG/d
ZJxne8g6HEPZNxzjASLk0wodJvmADssvr1vEKZNTzGeoksEi+NVfpDuucq7A/HQe3EvVR93NClVk
3MI36siMka4k1TFcEMuFsVXMQ7rm5TIZGGKDWArFhn4SSY0IYl1V7iUAPJy/KCe9Vr+LDSTwttLR
K61KxKt3LS93WjpUuTavlKEFcz8mmbkeVwgMjM/3YCAbAxc7kDiFQpN9hqKGt4k/wqQKapt4eAqP
oXUPNd67AaOeRIdNoMyH4y+4SY0g9l1x82+AzpDO/XZVVKWCnCcwQusk2mZjYiYhcroG0if69Kvm
wEphwDiyV/aY11MaPecMCQMbwnFiG6a1qablUaS+CnjG4q4Yc2X3iuSP7rIyOF7XJP2fJtuCICfq
kRw0U/gzQvZgMOjte1uFqC4F83Nwve+izTm26B3zBnYz+dv9FIN5OLXLj03yT+s8UtlvP2Z2ZnYj
2wO3YReYrjehEPE4E+TQDc3Ku1mqvhpWb1o0g/3rx7BSCVeDZNPBudAIAM2aaHBy0QayE394GjyK
SDKwwKopRq4AOTUYJOCPFkv2MnGhUjVebZ9TVWXQTGpdwRwYiPMZgL5IcDuCdNXw3G8XDf7xhzsy
i0LOwzy0lTAWfUKwcj16nXwvGZKppwSWRAuuZNQp2G4uEisNTV21KwNh41s4xT8Kb44FxoEpE1HH
ZBfrrwLwMUiM3e7mE9gSACWxaB5XGcUUIIOxcH37/Dw8Gaur1RXUps6Rd3AlWk72RjCglSduSSwQ
7ttjrixfaH1iJ/XuUt1UyL9M75NDzM+rSORBDM38zfhNQUs3Y7KOknzel+Cr/it0Y3OJWZNeTbm0
9VULA25O2/t/lgg1iLOrYyA5R7QPzmnammYuuOOlYgb5J3EGumkDHYMUnqq7roIzO9PNbXAhq8VX
BQCHoBi5zF7VoQq1Q+oEbkfmh7QXsG77S4sYTQJ6CglZ9AC6hQU40ZyGCMSkMfZqsAG/LXi165PY
NFa9FxUov9+01NuRuiV+gKfdDjK8rA4JwwV6tbbZmEGpZ4Gf9smnq3sPR3/tZPfO0FpwvzDr8HtK
B1jU6E9A5q4CaxPepereMolQGPaNxpF7K7yOPwo5iRpZgG5EnSeNKOsQFU71yGB50qLbnRoEerJf
PsSkD5HTcgphoqaezp/Qcz9R0hdh60PwmlMqnhL9H64P4ecUrVdCv52/H5FjFgGJ3o2DT9GsQZN4
D2NePBBSmAV+mxRRD9x6erapWMsL/H6zX4nAk9wWnQ+LQOu+g4A83DY4cYUnmWO2NGCUmFfOdvyX
l1NC3KaNCru8sRK2bBeV3U7K7vxb6QNc/vKIRdtlJ0rSDpAsP7MJDYcBpo7Wfu8fJ5AkufLjf2lK
7n6/scZmim0DeUc6H7HMXNEyU9gTa3S/mQCPW4G97ZOkBk+WZpzOGpwfabo+X391fPeOo3v4jGzJ
6ZiX0EOn5QDGZuHnhRJtaDWftHGS3vlzrPS0mms5G+UchkLeiQ27Hu324FLr6BsSMi7Z//4UngEE
aeap7LOgpQyRxPF449GJ7tYT04vqp+X3tH+MQgSLKzUsMj2ZfdyPeOFohB4mBN21zNUKxtyhCzZ8
q82dbdPz04cf5LB/6dRHi7aALp/9f2NZKhFFVOkuxZueFjo7kWwAppw+noJ+JjvbpFaMkl5yfUSQ
+/RGXz+lMRoQcoIz5UTnma0VcvdK+qLPMHRM+hX5D8Yi0BH5le3Lcy3DzUlOVe7eevfQQkFHblsp
ZsV8gSjF+2GtaY0FhlCx6JBuIdVAGCeg5rEVw0kXJyu9G/xV094o0UEiMOaREm6Y33A2vlhWBsTR
FjGOvzwnfkZu5P00dmsheZ62MSh8bi94FawbFKztyAeol/rfZtF7yJKENgWhePvhID0ZV/20rXtZ
JPfsf5seREvBPc75ldoAZ9buEdItxQjibT/LO8MMcMYhqfh1qYA2FKST0aOOM0oRQzPfS+5hF/Te
zVhDkdbNsmr9uQxVu40ZCUtLMKWu+MSSv2uxaVmYcFdHutt3inY3HDNnES9OguPK3OiFhjsA+B33
4V4b7PtgpZ5TXdXZ1DU0UmmfNJ0IMlOyax4h+1HA1bZK+FRTtdLZy/FV+DqLdswLbQWtlUUIKMu9
uMzQ0HAinyAVT2tGmvccNmZK//lP/oMXPKJ2/XzrXYp75A1s1QJdT3dM+eYMx/lyw9LpNHN39Hcx
iKQhq+nF4pX51DL7v83Izq5ZnAh/fuXzX806oSBjgpDkJ7dKUCjfNH65SS08aytnFlu9GVuvJqw+
UIhzNF5Dn30TnVs5s/KteWRWDRAmtRDiezRexjMZERUlpBzNPkxPPyfpXdvHOwvCC0uN+1ciHA4w
HxwnN8kMcQkYyxcuU1qmGMjJkbdwqFN8LmqrwTMG89DMU5tnscFik004SvSMwjV1t6CC+Riernls
+sybB79p9VPIvP15le4l3tYcWevey2QCYeEl36Sm/t/Fq5D6Sr+dXWdmzLXrD1BSqwKARsVG1j+l
0O/TQAGOefU+zqwVLuUQysf2VtSLpUqAvHkosnpkzis3HTOdwIXnORAUlVQeBpccZdZMLnVpvRwB
W1oLUWXMViDXkbEiJoXDi0SXIZ2wbO1bsv9AZOGQVHpRR1YYtGnNsw2lOR2tXwwZ8wsIbmkUWdOM
njMUE9scw81t/R3NRyJm1x1rCRM1bcXrHprn4r5gKunHv3SwG3ig06i8vZAUyIwY3YKr47MB/7GL
fTTChTyZwmGecyhW8+rgiNgvyxkDjWcLX2QhEXFOmZ26Atd3IK9EYd45Iwc6eca/Ryeo3xwt+0Mu
zv4F/tYZ0bMpYTwu5YPmv9VTDp8xpqBWOYieXyahQ21zf4xpZN9Ll3GTak0r7PbK608Trha7vw5y
t0jhUnerRdugrwlvLuXCjpyvqkYxjavmKoGiuTt2YdeHVs2ow5umBcZoAT8aTTUntErMuSRqd65i
MbJsSbL0M5FuWvKlaNVe7gXRDtFixpQtp/DHn9sdy7Qzk2rRhScL2DSSPg3jByPfm6hHEIoTD1rH
E63VH7zdaSlMCdV9hTsBS14yuTl0iUYCrjlJvA1tQMoAKsjQjqJQLQW+jAmSyQvq13KldRdpbKcX
Z4wbuA9OF8pYaQ0gNeziA+aiBzRMIx9bwX8SLJEKxxFL9KNA7Y6h9BHlp8zoF8M/Uvk1ENg4CufB
pPhIh1H5UQ5obFRn9H0JAqOzsuIrW4kncJvxIIH3wES9jqVzZwZ5TKRw8+Se1t9o03uHS+qASQ0s
rshJsxZr4RasBddZDmTC5oS6KlOz7uRShyEf0KDUUAd4ykzL+rufNh5hvRUh9nQF1w4gwK1pfp3Q
P6gJ6Hp3mqphOExfnfTwbKZYolrhXMeeel2BSG/oUXUaklkF/xsz252xTcSNdEYvYTPUwlvndpw4
Tg6i7L43fg/waNPuwvoDdgZXXI79ny5moB53ZUyUxSzAbJ2iEOnFXaXkJtCeCjroosPZExMtgppR
s4JMwR47fjVU2eWH42FF0346rHmrtF4+bfc2gI5ORGmG9U1JqmNzLl7wYOCJZBgWpW2sTYipZRlP
Rl6B++d9VXLY/hmNi3F+Rug7qodzOdunjIOPGohGMeNHcmm69vZyCEnl3GQcZPvhazww88jmKrv4
hX/IF97RoFgUJTnjMufoQ1vK4YJ3TggaWxjH1jq3pI89XysoxnAsFonHojgmTUBswBsYo1vZ+iBl
c1SbFiAwQQAYJpomR9cJE2/r52PW9K5lXAYDllKTqyQvn75045BSrQT0dJIaDNiCJD/VzYeVI+NO
SqUbQgBf3quM2CggZtvqnl/3jCPNKL2jGiTcQWZ3Znt4eFDf3xiZjXrP+XszgLxBVfaIK1R4pjAi
j4FJQrHIWSxVg6ntVP3VIjQELrXs+WVzc60bkMvfMW0Tzdwah8yMjiieJKRODXmGvK/wLKV19nuw
ODCU2zSsrOGk77elbtmVLQ3TJ7mB7BN3dw4wV2qmvstFnKEM62tjFSYy7Cp/cbF9VGaJC0x6Jk5M
NkIG/Qp5V5LBBEXHdwOYUiGLtfT/wY82drYDO8GHFqIJGCTeFf9E2Zw/mHIZpazMRRLUbG8iYMo8
Tp1PKvsrkiBGKzq7PQxx+eU8jA28JwROrpF980dgwFBduGZfGrUdjH76pJce8LQnieYZ2O7eD7Gg
MXHJ6FkKnUeKhW3U94oKFdQcxpv3pdeKEB9h9WVrCM/Ttks+SoyTpVX92hpcfg0QqZRtp6MNumyo
bwg8bApsuLlGhSJQDEk8XW84sH2kVf+Vofme3wfjeqh7MH2rAwQ+Zs7dR7WPzFQT7Xnr406KLZmF
Lxq09kuesMFIv+hxUMfTQ6k2OqHMoohsu8bMRnsaIZDXGHdA6xrme5hnAMEeXM5G7QBmB5vkclJN
oUcPfBfUXjjU3EIeSuiTo1UIkH9N7W8Bz7a41JRWcPH/TsprU4bn7+YCZn/Mx0caJyNbp+a0kLbq
wciCAoSX+ro699wS3EYwrHyTwj9MUO/uduILVWfWmxOoPUETZB+kpv1Pq6yfU6TPeLxa9uyWixgW
3LiaLddkSK/J2Pivzz/hB2r64KrEaVaj1zwtWfqZeIenkAIeI2OLEcypMCeTLIxiDLT4rtVqeJ9/
2+bDUONrjv+OLnCWLEUT3lG/1Q7+zuWuTg9BxrMm0WazXS6zw00bwjuuNlFbvYF2ls0b2aKDbOpK
m/fN63GwMifhpMowOZI8JSTafXkP75SXY3qGpFa0qkMR2kamVw+MqqQ9yDoGpKV/6+3zKwUBqTdx
QfRSUaSsqXL9f4oyU0vuHoTaSbuuHX8gQx9vhNzFSDaQEu6u9yYQQ7L8mgo2AfcXW4+BvE6MxdMn
gzDm0ocxcmJt+sULQuf6uyQ5up4XIeXVF1gqZYJMxhYjhju8Rx0Z90qYY7p+k2pRL5Uxli0oIfec
79mjRv3fYkXBvA+OBLCNPTvXm2WHkyoT+fW55O0phFvXZ85H11EbcZr5+bnq2rjnMqeEdnYri3q/
5DlcNCSxWUWKL8j1YoP/Sslb1GfRGT+Vfnq6SX0RdsfY1Q+aH9kjbwYTUOH1ceLgG2wLUNIgSBzX
N403mtip97pEd60wry1Ib87ee/SfhlQDP4e4IfV1hs2OiF62T0io7KgY8CmMBapAzIxqZ8DIStBz
PEqHTpWE7aGm60audin4XnUorS6kwCbnocb2UyJbkOd5/B+rTh9aThy0otseo6APSuZxHQELxsGx
krIUC4eQxfQiEeWg5zKwPVFa/deth7x8mPLbqEXuPCC/EcnQt/d248WC30stRxixfm+brCMTaNkX
hfoqZnDHMoYiMHx/z/z/eBnnU8aEubNA0fo3fYFjpBgFwvRS6Gzv21uLirEHhBSq1tnqXnu4OP8S
Z1k5Te5BX+hjpO9HQS1CmIYpJXOZgkJLxJcbW7GQw0C2Dl3A5LxbPGOXhX/CK9p3uKJt8eaFdGAY
JzPuw61flyo7sGBIeRC7I6NQsEVulRB3XqD88fAtglotZytXnOLkKKThlcn8ZDDJBvs13DfZnicI
WNfj7ASt9GIizwrp7qKm03ThpralVYi9VKB1W3IchQhCOdFD6WDk48IHgmLfi02a+f+qSrJ2zqgL
4dsLLNGlrVWEsQ1irkI0jJRGrepbc9xAZMdNpZ5262fFxId6u+Fbs7wB3qBXjgI8Wr/E4UTXXXWb
QqMVEIo0oMlXu9730LJIpwVUPZfwqNArJhOjvvev4k8A9QDj+BKCsVCgOwqZ99I8lsI9SCvuabro
k868cH3nNm7d09qxRagvo//xDQMQHfrUBlaQtX55UhA/HQ5gd2Bx64DocC4vkDjctIRmc0L1W4hq
DPCa02bJ9kYL+SyNN75s4gKGIEE2z2RIt7CylxR5fPM3+SKcngUVUfYxtAuarYFEYMwqRpbPF85l
JkA3TSxGh1TztL/JLI3Gfomcse4wcfVi7cComkDjOvK9Sf5K0ElcxfH7oCKi/ARLGBfNHQ181mbo
A2uDtXGmWAiaUVhgzJmvqDRvGCh9iyJG28PLtJFnQLsCT40OUyFPqPZ0iVkfivwgRkbDPr0qxNda
IUarLsnqDuFUGesdnQ4/kpOsg+e6j6A2nWS3SeKUYcNcVb+uCwTerNT4pFKbDk8xIZ5d23dqx02z
rPKCXob7ggl0CoEl5QEiFgvghrObPT7ceWXjuEXMWd3GWUIH680ROT+DcNh4kbkj4eDAVyzNk+8T
pjlLmdV53Zn34FbVc40sxUE5FH2hr6/xbQ38LARUQKGhrAyQ17Ml4Sg7PL/jHTXwNn6Vsofj6vsH
TVEOsI4Nk4UUDEjgn0SwnMqYAkZjvAhROEBrF3Oqix1EY7yQNDYZjjk368jrus5ZujknHevB4dWq
tvDbS7BeCl2T227aSgHCxG8fpz0BmhhfXszQkFTqDJOj+pPBlM4JCvkjpk8c5bMXjvXZluAx7HOv
HCTtlvcI7rWlzhqpPUas1Pld0Tcm4vK/4GlZT4mr3Uub5RYmgow8TXJafQ4zgjHe0HhBfqhZM8zT
Vocylxx7wV/M9hSZhkPbdCD+VE4CNNdBFNAK/WZDLZoZJQkbg+jE1RIX66HBmP8IUsKzBXKsJjX5
Dd5KXBAe6DzkglkG79Zz5TQhYkPsEmH7QfBduZiS0vJgrRbUgyxX0fUMbdBtqvV24bnVf0gBhN9c
dSKxA+rzQ9MGQVmzSkWGfQG3RjaRnOykjUBsCDYEs4dpcp00o+XCDlnuTSnPk+sbwcZtbSN9bbO8
1R9j1KL4hJqnGBqh7BcHK2FR0NZIKCzKFaW8h9/oAWcZVPn+AJDBTEp1rzTicCGy72SaVrgYu6QT
S/KFtlXa/WIyyWUV3h/9Ue0LJoO6qQAFIEp5Hk2obNG5yq5D4vQHObtxFaFvlMETzV9ba8Nsqeyj
zaSMSJkM7+rve7ltlwclMe3t3v1RORy1aPotA4Q3ake4Z6T4K/4jzGyYculgpAzwtVqo49LS/yUp
dCI+iHwqzlggfQJjz41yOX8ylzyxLcPpQ0NswvjoDGhwrbLNW2NiXSCbaiF69l2KUswlUaAxmTuU
LAM06luS9fCfV+xtJQ/piLQcRUjnYVHigZv2hAAYJEBMsQkFuDRdcQC35/DXPLv9RxZkJ0nop9zR
uzkGbsr40KWsRhSAxuECTifD7TB5qpwvi8n9riU/l4DvEdGR+sdQgdKw/hB/QXYTi9fTuNcav2d6
HppCNPhXO9DpWyoFbqzqfnYS0O/jEto67E16OoaSzdqKvimHurAdCvVbIOvpHNRoS97AbQptc7Vu
p3FYmO775yyF73JRVLwXyt/ZXoNQS3VMLdKTsKNJWXus8mJ13ikFq/72NnId9M3B/L2ids+obH+6
bJ9jTyGcRZRo9M5FIANoGxjbJtwZmnMF3pLNdIAbWMArGG3v7yUhm8xz18fle1jlWRIZG+aklPS9
GLeBhlbrskqojFf9cXNSyllqWHvo+9hMNXCzy6X2bkcQRebtpxs6xzVHOqgczwwrN2FTpniH0Gyp
lvA2cJnOXEQRlNl/ATy20sFaRaY2ifsj/UZ1wmFLR/vG6u47njuuX6+jYE9NCPFwoPSBR2fcPCPy
lYijB/FlNJ8WJtbUjJPgD4C8lh0N+Wmi0HpwHnHqFdPFHrOEyPvIIZ4r1s0mXWkhlduIMUhmSf1W
6uLtGL3cFD0G8VFX47HHfNhARCVNrc8j4gh+VvsZCu4OV2AbtpfzAPLH4759lNeaRtfgAh/9KW99
aabrn7hncvdIO4HgvpUYKYexXZHv7kDjxPQFW91r47/pZh+q6fN9wWYXj/2AXfDdgPdN241bzrE1
vbbe6WKTfKE8xTMpjgYGIEXBLULcpd9KKXyIqC58WZ0vP3b4sAIOUaqFDCiijiimFOC8Hl50NDA/
LUcq5vf33JvT8cWfnP/DGi27H8JPIpjtZQJehPUPMMliJnvNrFsYZc/Gh2OaHffN9TfUxtYZunot
EF1dRFV366TJZAQZHI0wKXQ8+Wr517IyUFcDUbmOBJceA3G1V0wnQfckGWxsIvIItGeW7nY9Eb1j
JSd6k1IZkVVeaqckZvx8KZZsrzQJtaxVhpyHAIFHaHXO8OSCMvzzXNwx420abSUvxcR0CuBJiICV
g1Q6zY+QmK1KM91ZozBAiWt0L0h98LZ5tgLYHiszQm6/qfBgEyUqDS3PTFsjsCApYRHHO3opwAqO
gmkYYny6GS+84MQlxAZDb41tCx/Jn+H7fbj+IBa2mmYw4bqy+WpKEhgOZVIlJS9D+h3uMDFC7+sR
LVHCyMYQI2F7R7t2wus8i5gCN8a5bnxtCTCOotlHQgiKIC3o5Gtd7S4kAQ6/ye/RvJ95ij4Ug6x5
aRW/BrP/DZnnjkSLd3Oqh2FtbVS89odRh4y+SeAKmbL4sgKTkuIBWvi6cKG9hB6Rw7gTYGDp7pyh
U+7xk+oeCLhhFGjKXbpepetCoY58Ksjaa9oih7mlST93UYMsJGSxFf7TOUfNxi5g63yHn+9rdVsV
ripEhAQ3PPlX14q1fiZcsuOprG5PkJufdSxPkjV9uahgiNBBQYQYbt7r34pjsVy0Opu/bU4+ZdCT
g14UaYa9tj2/0A4sOdHbZqWCZNucZRyHY9K/MY5r7yJojKhAxIUnfuRWd4UrQvIYKMPHIT5atCuK
W8RZlcvzLd1hcwejH5dFdfOHNu+3Q+z6uG58QHprnPpGSOXlNvn+kL6fsqYyVZ63IpmGfAUCMpv4
F/JSREvsuJ5ht9bUbowtuEJ0tcGP313xbyIjNDTewI2Y2PQOS3P1uC77QAnPAMzhTDMwPMuTcV6x
o3VkZS6OzLZxzNDHD1hcrRU/eRiqOxJvcJBO3ZD0GjcKIJmh6JG2Ckn711ovGTTiuJHO+mSGlR3Q
AujKMLPE9hdohT0jrMRxlj/zwKjvoR+ycpkXK/tHFmO/EIB+TSV9a/2KuCCcCbKlK44rWKdQEpFs
8VJ8ZT/CQo9bY8kYzOrv3hGD8n2yeHejUKxtl9eGlm9tDw9CC7dFcjdEFXLlYC+0jovkkHMjfRNG
bXWffyslseJqjndfQ+W/ZGQt+JMZcCh47ZoXwWps50GQ1tMotkegb5vMAo3jhKH1ZYDYkk9U0/s+
HpWIG3smPHbkZSZjXVnnUua8ap9lJSjzcWaIogXZGfj1+nhN3IUF4pS0B2D8kpMse3U3nUAaGXev
qXdhkwdodOebNPbvcR1VXJyCiVwEB0PEjvKi33M8XgfQPYZbwKs8bIVAFE6D7XfWy8MLmVCNkXoU
qoVdbRfYdT4HGMzdUb3PE+jz4JwVCR6yqM9Hho2mTpYCfLsA9zo1OTPewsSXqKH2002FXvm8E+7g
pilEcXijBFoN7uxqWBbo7AXjczmcWBS7X30pcQ1n4IjbfbUhYoXb5fJJOoWqE+PiWtBjwJa9TTAi
x+z5sCEiZSt4ltQsRXd53/jl0zePCnPPddZ9fYskfi6RlFCCAXQF3YpaX2ebvO7WgaK31T71KMhD
wPEkTMmEp2KoDJjaHi5mpeL38Wq2IoYy/wlpH75rHpVp3dcfAP27roh70DEm0WGAhmW9dd/hxymz
F1pljDVmUip8tn8FuhfJLWapU6WByNbs6wdkrDIfWMh5zRRCuwdc/znHnxX7on1YHfH7aYhX55Z1
5kysv1lrUKZTlVN0z8+GSD4JwqeYW6s+Ts7nctJJTaPiX2aOU+A4Zkps3ZnU6LeFV/hKRGrBIWnc
/yZ1ZLSF4USZVE602KkEIhooxtimPmPqs55vHSO277UeIyyKYLlNrNzFYeiA3WPf7MA3kXWnweXW
z+PiF1b1aCLKWZNyd7Lf8AcYyJGg1QSFIXxpe4ORPWNaaMCB8v+owTLEOnxSG+B5brgSmOwlLIV9
7gX3G65cgwaPgxhRloCKuDtVbgAOxRtzZbt9pMBTIIro2gQ2NnSsAWysYy7jYDEY2t/vqqD/DMCS
bhU+S/yR63iDT8cAckrWfypf2UltjPM+9HnB32dbOr2KeQcGlK8dyKDnGzyPykSZ02tiCWC0HXGH
wwEJLGoFOsNjBWrPGCbRVicwoZ+zFMSGN5rfYz+X0KltmUHztzVBLpAYkylMM7E8HTy/xaCm/pUC
rWEdf8lVlOpeqKrCH10nVI75mJNWBVS0Ap2z2ZVmY/MoN9ibD6B3wVGqhwgQV4QYqytGqlWuU2wu
3jt7ifNapAvawY5msyXjXCjqNYGReUtGJBUQZ8/1k+gg1fbwS3zwZCMooqr0SQY3+XkMT1ARs0c8
7QWTbVWByEhSin4VAU9iHjJ5BgBR7UQVJL3B1ehg5xNlvS5pmd/rZeuLKjSIBvh864wcBzb+6M4Z
U7+uCsrqEDTBYvbdjGPWs3ufH/9pJj0bTYmGkhzQBCWm7Ex6yLTrPoTFkUXyWipD8i8xkO/dCkmf
Bx/1zFCwLdjLRhQEgvTdYmz1gEomLOga2lWGCJsIXyFXEu0VXPeF7rByVQi3K1bAepVwmTRZ5vQd
KPYASNiuKV0ZoLqsxrp7hSMI86IQkZ7aUSNk89ci2iawLDSZLuaZzMn5R+QHkzpEb+DSjl0IZZob
hJA1zsMIASwRV7wZyIPm8IPl9mMBH17L2PJ49S1lGjSnfrh0frGpjXan/5k3hwEP1vOv2VDYVqaC
ByEj0HbYBI8ubSHXoz1fx8Sd5IGZByD6JKxomIT8aCylu6zKFOU0Cwx4WGCX4iaXUhPA7QOXIst8
uTl/lQsYXrDVg5UXjt41DViI6IF6/zJpbxIQ3qx5KB0ninO30X62xRLVG8cvtzlR6xeQiuko6fEj
INlw89vTs4vhvGp8sAWh3vPURPEwKLgIhm8gawirkKc9pp3syi3d4Yy5+NDB3zO6j+vCFBYp3tAZ
PuGIkdhn1yx9hkugwA1eqtzj1Qq2nwUjuff8aaL8G8ZgD423kBQkcGJGPXC62vu6g+PnHUU6BLhp
pNJvrQVbRjZLBPTFEN6H6uWstnAXVzyKOcwDXlvAYo7ZeKkdyLdmrXaPhw2wuDx9izvfXSwUSQr1
avzEvaNtNuilZS1BoAKLqgjpNPqW5wR9WDv7zEz1NLhIsbeO090rtb1g3M49ohBcAuhyvbgurmGA
u9e+Z0JVZxHaKQAr47LyouV9OTMH/HhJvomxSKTB/ZdGP07WCQQ6dFTjRO2x0qalYs2bQ3yaDzu5
8X+Ci18kUN4jrgHbko79ABndOZ9W6cFsZF4xg8o2/cQ80UWgAmdr5V0cztTYig15Ml/Y3o2cnSPW
9oYCiBYrLc2ZRU/ARLe0KRTDO4g/TiaotUsGEBBU5gLIaLPoIq5PAcOpTMHDk9Hf2Wu0Ki7RVpuJ
qZ9+Rqf7chV4YYHcSPGHHgy18TTNAyi10iWxmYjQDtubmNW15oGE4A+DnknxSmzlSOxvGZi301nM
CBVLOMoFgeQ2NcXBhmM3+9SII4xQCzX6ZJxjxneHl9eYoy+STeu5AiYpkNGLj2fB7GInjAzXhemz
O94IrfW4U7hHHk91AzY9dyUkyYNn0S+SWtM/xIOgM1KWia5YR71fZhBWdcV6hV3vGgyzcVfDv89B
KAFHSIXascm/iKAcScADmvbccCTgKvXPExZgjm0SIwQKk5Hpsc3ZIAN1hPWoONDCZqJlXalKF4uc
qPu7/nbuVme1bt4be1ATxyXAIEgfW6cGRFa61MT0frlIfc+haC7arIQEUwvJncO2GZTHSy08N3wf
vDGK4xS4P0Gw0UyRppbOOh8migjhT//MO6qqJXp8RkfWlH4NL/X+FQrvCFGNX6D5wiiRJibDQCum
2EjCHKMrgZ0xxRLO5/JmE1KshgEjoiAFrycPUKGuWEhmVGgDqbf37DY2JCbxAJbAez39Tfmn1vvz
l/+ZxzSkXxQ/nnv6cEe0VyFHTrNNKNgHx9qe7eTLklAyTpGSDgbovSQSTfbBWifImuB3d6iwq6yZ
FyCT1pJsp5ATB1t3Aa7y/rjalM7eq4e8nA8zrOpr1hZXiGZdx77dz5PYPt5ISkZPUb768ynZF/Yd
NdBU9frHFQplD5Xz+3FGuPWLwnPRX4/0Ih5fLQHnSPnZCdsizwTq04F9hkNxFATjm+CqV6QU/993
7dzgFewB6gJPZq3Dbl0SEVDCQ0lTO5HZENpeVhhNmHCG9kWBNnQfAeaxTCwNlQfSWFKk0Hi5xR9u
GqqJgkqIOGzCjhfsC1JiWzViJ3392UOiXS5fDae3EsP6f453mcttK3I8SrDf5YM+cxRWxRgAhP5Q
6nCA0f3cc4/LbBFvbLRn85W7/kOoTvdySuSxX8pVfyRcId/lmzJ0S+AJPHgXcMXUWJpduU1X1BT7
UVdEu8EanTfmgHtCZOgHxyTTwgy5m5GgnR5ybvSbwg/IiFG6bMnNXNcNdWum9SnAoRqPJbUYQd8/
CJRap3xLlqb/lY2xkSMdctzG47ZcYYm6/HeP7BckpsN4EpvE2wk1XIpqWDUPJ5expSpY+suS7hFH
RDe+dH2mbssh7+sauGKhb8BzVldNl70M8ai9/4IHh1U/lBLET520iKyjOQNuInwfM+MYglKwM1C1
S71cVx+fhxb+81hUsBSAZU6dfzqAlXHaD5ZZYWvJ4ZJ9HmGX5aBlkeuQCnzIfQgtWpynL7Q67f3N
GZIaZxStbxwsenz5pWUZK1WGhQDUzKnqwV2ka8RwamdOHSmBRN3L+z1PuDWPBpZEB1qL0DZoOgGp
kcym+HtXI8/LrKLIbxTS51ImY0iNuHj/8fa1xTAfMvD/k9V5yTdaDaNi9XmIBl4eJnFjpiPK2dq3
PMOhHJyNTzJ/ZoglmXHjPprffOEcwSfWazOPoTCp58uBwZeE76AtcD1A7bNO8AC0paMdxiiaYlwB
ifmp0ySqGbi5SpNwUNRfGO353m4P896D2ekRjgNj3bdTGqojfAlEswEUePwRClSh2MEMDlbNnmoE
lAfaWEKUj1RTD/mfu+0WRR6P2lyMz0fPl/VXn7r4E2VxulUxs+rJTn6l3Xb3xIN/EhpJkbWwpik1
VQU7+BWKGX8TZzrPPKfISWWFub8DgRtAEQPPdBoneKQd+ssKTpFQi4Y+S+Yjc863R4U83zQGiHET
Ke8Byakb9MavmQpWMxPq3R2UQq7tDWPTZTyXe0dR5ESjdNw5OzE7/FGgGmM5iO/wl/6t+9JKhGcL
wctc5IS4/MwLtLzIBWmGiB1i6RLWv9WlTty3HaZvMaTF3LLMcxaaNn3tvTFYw9hhHsN5QRP4HChg
9D21LiMfvJ+qlnZLU0fZzXCnbpno+vD1aUsnrXLi9tb3jXfYm0T2yGQsEF24uEHhnVPEJzPfOe7X
tkaoDd6LiBM92p1qkm/VNoMGF6g6InvUcE0Ived3DFPMaLRUbFAuqOKUHwcRY66oCCgJk8HCqdAI
WQEPaUQMBlKqxKmZr8gKfksRirJ73EcWIOekQMsDWdVkhQGF+ZDoZNuwc512NgoDPWcnJ5xjwaZ/
yjwl2fn75bhv//pwKJCSWG3C/CNUzGj8nKQuTEqy0OAqoeSdT7ISWkTXCjwqSH1aew9VZ33xwizz
H6tPi5dSHd5ls2pKdnLkqLDBT2MRAmBJ6NGOhVGNNzjoo+v/ewLbRbKMmnGsosvgz9nirefIcrG6
xPKCNE0FRMMGNepnqcs+TFXuTvRGeFVeiBO1c+LisGHOWIPAeFl8IiwaENzrNdQ+h7vcBRyg8wNB
4AEZCZwShgXhZrJ3rLF8iviGCFaiPfGMTXdazGJi2J4w8Ny/HIM8qhT7Yrl27AdYIu3GeRka8ZBh
u2Cev9eLGwiDmZkeQUXiuLuPMcAf3bZZRRjKhz7WwOds1mPTI6ZJeb8ulMOYMm/7GIJuPDSMaRy3
EqMISuzAitzGmC550hoeB76PRcVusEofftWd6pUREvn/QH1qhotSYw/ZtB1R9FVwJgiVcCXVjV5+
naaeRdyrtEfXB0BlOJH259z1aZEMFFZ9ahJH6vP3hOJVC11Dk8RlrtYCJIva/os+rDzIUFEMlPBp
y0RF6R0iymHWDmmDhOux8hRL6Hb+HaMgAVXpWCuA+iFgJoeUlSDgJ6rMx6als6K8uX8wYqR6yv2g
3PFtwhVQOXPoKi9aYTPfqamo5sFcvfa6flXL2+LAe8lrFWSXrhqHkRjQETjzCj+bL4opOM1DB5mD
bcptv+hFrIFBFBsZp5K2PVLamMBpRcdjTzx2tJzZAhAGUUTSpaPiV+EXhXvGw4BNadWlTHA5n0OW
fk+mye7mNEoZrv+aEb0QKQW3vHkvMU+xDY1CH+cuftgeNQk+zxQeY1bGsl8JEe5i/uKsTW0URu89
QDdqdmLXhItTxN3QG4ZOawDg7ctyuSrt+RhK9LFXQ05LeOa7FV6Q2lvomq8r8063q7kw8U6rTRMJ
zfVetYZ+B4rHBkdLw3B8miwK0Nrb2KYiWn9Zts9RRevrDVomgWEicLsHcpU1x2OeDI5iH+3RuKeo
WdH1gMaJxVziCGV3mxRu/8Ph3CiGiGMK7M/fA3KJu4wDPjn3hnB1xvbWuq79voED6uvOyd9NRe93
WQlC1ySFS4z2bg74w0Ikvnf0TfljM/AZlWAmUFBuKE1PQYO01zBRDuC0P6SwdolK2779ptvx/YFU
EfucunGaf4ojM05rSbDOeJSJON/j2iwpXNK2elb/dzz9PB72IZth9au8b2Ppz2d0GIsWODP5A166
+CghRMYykf3+dVeNpukzEFR5rR2cwq8G01Q2qrMEYcCjJyxe3imivtcBV7NdneMUwEepbyqCGflF
Ottcew1C8V7HN3Ul8kYDUyhztTs0q8xNYLfz4gOTJSK6Fw/BQTqeuinwOrbXxzjV+ng3muRyh6yy
HCwqKC3cWhhKsr/g5NjfW3Mlk78Qw0EC8MN38y66iOukQ7yTE7xsKsTH9dGwU1NsDXOSgbJ5f1xI
0QirsVegVle9SRCGRwdPx5xHW8DwuHgWx+dPiCVuZq3ttVhAT0qnVPXevl49bzN7WWEhfreORDuh
LR1hbZTmWesHE8pbUJineIY3wAjBjMWtXZ7tY3VGC1VGIAEkdkZ31KcEvzgyVeqPrfxmOREjj1xW
jkoWUsN14bpnM+tnQfSGgBfVl5v77b1m1skZ/He05wKcfe0QLaSZ+eHMfUDmG5Uj35jvigTn6QYD
U6HltSkZKBAkk7Ld5hRBOB+mx9WkDxyKh5Vwl+9M7zNo9g2kmdzJFx4cQ6epYJ24G2cjuN5cvCRY
O0Mf9ZzewNfeeCArW4AiXRNHL1+bYcfpXNmFEe6WpA0m07Q6hDlsJTTHCX3Z30HDyHVTy0Ec+OqK
FcOprahMZhDpumE87uQKngn1J5QWYO2ef7AdgcLhnEw7jnWCMsq3EDL5b1qHTvxXL952DURkvWQs
Ifh/wkCtkqFE57ydZRYEQolMzfbwlDP/P70wizrxUQxl93V5ZSEUyF1s+y4lUBgpnMmGYDd6ATb3
8TEJ+rh8/7C4whOQirVBFyAxPGIVpZzvvfIwfj3mBtXc1HetIbPfiaDdHMvg0mD6TXhqj07zHZn4
7aZXYHWhpCGh103IpXDfXYSs972SN493hhd5RnaLd7ccPYJDE/7NFXNnvOBfy8cFSHSrm147P7Ir
IDlHzwiqVoAWHCiiMaFh+qWyGBkPbXoDh1Jk8hH5FR5IXrcxoRkhgZIcIdwfr1lJ5593daYUgIpq
mGz1FWvESeKsnBK7XkB8x/sfW8+cZbPenpu8ypXOsmlNF+cYusGVMGrXSOa2I0+TrR78wgDjJ65v
gErYRo6UiwRuX2HYlOfOh8uu+gWP7ouXalcYLizZo+NJSsyGb+SzMLyKt6WUg5CXH4afQxDBZgA/
+waH4+OtsiMPjQIvAj1vJgu0WmwXRFZeJObdHhJkrw1Ss28gAUvfQsVxincNaWuOUh+RfQIATZ//
/tNkekB0Wxa7aShaNbz4FbfIKbv45jIxy+ndT+HtVFprUrZJkCTJgXOkQ0GekaKxd4AUc8UC6Kak
mLyJ5LotIyM2MsfNzZWIULbME7PMU3BgB0tjvF/PPi6kpI/+ztRmGjByFguqatg1ED8r11pohdzI
PVxy1wSmUBNuCjBu8AbdwEJopUVHJ2AnWB7ujGe3n5WUwlrGpOJ1ayDOB71AWu7WQ5Hzs8ifrh/0
nCjdKk73gT/16AuscGiBxvV072iKA0lqdnRib/FaucOAYY/3fjj8mkJhSiM7/hFgEizpj03D9VBJ
2mQEiYM1WlTXcqajy4nDowl9uWOQdFeBTBePsr/y5FqnFpfZatqWGWI+DWnWBWNtPpayDJlD5AK+
7xQiaXzReFtBXNxRLzHlHwe+jVY7/z8rAm9IfNUpZvNPydGgfZGK0aCP0phQq48T8OBqLMnBpTWn
twCqayPpI9EUdcIkL3WgUQ29ih87i5O7wWEuxsA16rtaBuhw1LI6zzomxIG8Y9NEyybfSs+e154P
DU5KDo0vbHgVCvBAnsvGFsDIYccXu+RPtJyBmh+pqLyVPCe7aZGt8gGzvv4ZFBok2uv2r/VUZQs5
AlPc6kp9xSmBUuKeke8Ymb3ETVeNtU5xCg/WvmQhgAgWLcajaYcyQwkwCCcYshce/DyOnkPrW6y0
uie6wcpbAdu5gkLM9JeEj0jzsE/P9g2Bn+emdwWZtVwkoFfk6jABjzfIN6Ol/tiOw2ONdvoXfwSB
CygaHYpmupgllP70lvh8lJMAh3J93OJGJYYVgveNookejz0jLQRq/EFKF64sa402C7P7bJh/VcQD
6cr5xmAl4XDyQqciOVYHHxYStpoNtMUatkL880yd0oI2f56d4pSDnQJA9LiP1IunwlIalSHoZOAs
snb7fma+zGexvPR6F56vaPBh6SuN6v/y+Hiiiu9LsQOlUY/M2xmnLsT0QLwkET0qgqyKU3jK5GdH
GWmS7CcYsbzgV7BSc2+WCNGUEnYZJ9g79PSrHA1ris0Znkgtdi2EDS48n3d8/kMmPbaTrts6twLh
km0Pcu25aDFlREtcT9N3mQljrRsJiL2go5CfIPrBx7ckX3QRRjYPB0Nu8f5jvRR3RDLePclFD3xL
FIVnhfxBKsJbQ00fHm0BnfIGXy8PR7ymhjqccRDicG001VRncFNcehLdMatEF0f8YIH5J/FwLkcx
4STAIr3y1lpVW87zE39+eg3xBML7TMXN+Zsr420rhUrwJBpPIEC4xcBTK862N9mUJs0s0WM/oZkk
zqIyQirTauGB0657Xh9OR4CLFxliig4U8m6KjR4SQ98GQRbU9oeH3eOJEQXL6HQ7tD0YXGRsxW9Q
ZKwcySxv+RKoDNIsiTOkYbuFoqQrGJ00hD3/eUmwCWZp79kuTVcxtVW6KplWv35LHAs4hRIgKMRO
EUtXqZN1qhp7hB0VpjCfmM2lEir7/MUN2D7ILiBWDpsHrz5JpE570hSjKtV+MvUTHxcFh3/P7M6D
qAKUayC6Ak+2+tnXKkmo3YL1brha8+tdRKOrhzcUMrFMgYMDQCJroxukbglGR+ywvN52nPFCv1Q/
7/aKpPpv/vityvvbnGHhPyCWz+pddJHg+kQqMvZfXyhfvyHNqzTt0KXFS/iN4Crdip8hgbNtEVp6
kOd993Mn8E6kLTND7lDB+7FQg5m/eBGpXxxIzi3aZbmngBwJwAfJjiTIVrs7XMQ1ANetBzDdT6jB
OORbbKEjpEwV6SoN0+Mdmd7coOZpPIGJxmcOPGg4ad7KQfVBPcJxXpiw6PfOIUFVQYgw7eyY9I8d
89d01zGJzz0tfqZZHpVJXaaU657dOPJ8zkC9LDg+CMjaDcG/aqodhR43oGpSlFWYNalksinL0pbP
+V6ulCFyPGoPwyVD9ZrWiRFqahjCBoTaa5yGcxcG9dbDAH0PucNxcW65MoTGeKPnWhVBqw6cQFRm
rVjYRZDCTTBBIriCIGaE8acBrV8i514Xe0rasto0at+L+avSvYtnylyRIUF/6JY6cpPkQIBI2kZx
MHSkiMfLzF7PcRLlpXYxbRvfXk09QKHqEgbogAt8sggyhwBq/LVEZAZvrp5xqUUZP5DvhMO8zjrE
2mDfurPSIpTyvdOVC1GaoKK6ECGAu52jruTT/TYfZEBkINo0uZ7YuGUX3YQBiU4X27xyclM9ctj8
tFF1iNige39l6fxaWYcCbgxsr+KrxvRoCi/s6aklS2uxPB3ks2F6M0AShy6gk16FJBAuHPx6YO1d
k6TMsfcrwS4BZQol2FtC2wO8KJ821hWGX88Gpp6caXGneSzHflt2NUpdS9PEbBe46h+ouRfKR0pA
Nld2lLv+pYN7tLBvkUVM3sqnZfl7NfErCGCbGE9b0LNRRImcOjySvEvCle45RTPL5v9vLQuADmP0
/NO+IIVDZpeIyyF98oQQ5fvY/RZhWj2vH3uiHpjjskrlcmIVj07gnjwvjmxS03tZ+PdY7LxR+nzA
DTLdFUQstX1nyRSBSMYiwcQgNjZ7cODfIoxMEnZOhiEH0wDL6wFt/fBpMeDLq3huPnR8CuAP8f1U
pYPdro0B5C/Zc5QJFy7uIFNMonthrGtSuovBh2Fc0gPjL3szo6FdweqLL9Y9BbogPhUZLpWmb5qb
Tu1Lx4bHsY77zFKmR9GMLdDBabn036cjyjXVQiXAOPkXkUMQ5hMP9W8nkam3eP4bPuTNypeqi4gh
W6qz+lBUjP2WYtWgyMu7lu/NJKDdBX1f2Kq0SRnALhcIj9om06UqRqowRmkCze0ie3Wh4I0yec2m
tIPLhNyfUqon0xg+cYsJR30cR/g7F65DT0B464wvX6C3DDTPbDYJilci9X8LjpNfAHI57+8oTsnh
XqJqqiu0rDfihUxasMiuU7eJNvK5+u2vtB2kUQJBZeuzu7WSldupZLad5TDyA7YbFLlrqIyXYcwX
x2m5iysAZnrylJVNb+ZRnsS76tJoVgXVYqYr++tdpS+pmrAE1UWstPvp2JF/ycD6fdOLdtVX7S1n
Ue3wxI/tquPTa/Ws4tOoIxz0UOAvPN2WCseUEavl4dksPLCZOvXgyOqWGoPybsMNYgmI8oGNupfi
5WnynQEVbsfr4z0WJ2vz1bw0s3q3ECmu27e0ixpPuEZ7C1krIs9hqgAz9nJlLH978eTz3cDkg8se
xVRevlaZqUrqJSqT5FCuBlvFBdqIpmH7IXSbueXWRIHVozBy79ktyUCERco1S+5xFRCy1EbE7i39
GlevsaNvloRmsHSuleWfyQdlcsYjwK5reMKBV67fjQmkaDw5fy5Wr/xI9zdO9fzevSIT9k0TUdxw
Wi+UFYDL4ey9XyvkuxvPice+wjdqzFW1aOd26wu2I8BqFeFWkMIY5HktlnrzXf4xjvMEEShjVYvH
O8w9Kfa4Bf5Uf2IHy7sQ4FIO/7INXg+6Uj+lZAvqaZhr6+u53Q4P9yJ6mQTW0UYEYBn38vKMx1QA
3uJCxJA6bM/n4Pdz6v4SaRHOhW3ZqnRfdkzhcWO+jze/ehTvEdHV+ICyiE1S9a7jT+2CierZTZoU
3v0LrOc4HBRaboGk1zuYMuRp8MjVwDMYG8+kw+FwkjZiLOwfHoUaAO7L481As0c47rYgT8vP+VS8
X/opBAqrx2mOLe2E/SitpXVpgTuQbO5QyvQb7GIrAFe4ZzJdPgBT+3Ig6HsjC5YiieDrPMAJVRr3
F/1WhKw65PBZTHb1Mppmet8RkMzPdUuxnuXO51R/zf2Qw6xQIrT+UkerG8Er4oQ09sRO2lhGo7HX
lw9UWBazVfrFX+aq5FRHNRQV9+vmiFdh+j4KMnLGJZS/WYPBpwVwf7ga7K8tGV+P1JVUgDy5CLsy
1FZ2SRpFBMIOYx+R7DPBTtU1M2FpJIO5PXDWjkp13j69J8Hk/0DIh/Q6Bo9Uc2sgD9SdOHBWPEvb
JSQFjEq67P/8ZJv2hYANN1KEtFWa/BwqRLHnM1geZFDxsuJtoDVA8VlkqdGnIi9u1AuN9eGqYWsP
Hy8otf66e8JKi3qdImTWrXEjt4w9CgfwnUaFWMQUQ+HbRCNW8bg84TIHd3+s7Gkz7KFbu5FbLy/I
Mzb+IJsqcxrK1SuvtEPIIrIC04D+JlJO9ZphD/9/fLSmMHL2q+Zu8vogpyN5HpzbY76YMBruTspR
83UfP2C0kkWfWr3lys+4f/3AukX//WQrBDV/dT39xe2kpxLKsloTgC3QOAReGyK6ln+Rs9gkWdsa
SpUOB5MIML8AtwidrguyE7isHXqSqyxNkPqNcwwyNmpfTwrFnNl2BHkMKBoLHvXmnKl+bgi9dOEG
r3J9lM/WkshUCN9bolNu989OeBQWKQjTGxCzhE6c8W4KGI8xjTGCM+YcnTkbrqKxfSVTss0KR9hQ
p9X8Pu/y5PV9TxSlc1ao3SRxCk1CjQkBjJ+z7d9cKz+tgwqMSZb8IXa67PswnxAfdJnDQPqNQn7B
dyXsbcAOqw+0rS9lMxRJfA4C7G3HHy0w8NKtPfGD4caJP/9mR+Kd4bXR/+N4b6FWU2QR9EMq8VUJ
jahxR+d7WXTYgGzozN9+932GhmJBSDq9p5bQMqO7d39odgPFqzEDU6hOxohLn/l/0y8/qX0qBbyL
+4x5NU6IAtYAUR6H3ewG/F/snTLJfkBecoSaTkJ7uXViPyMtjpwc7fsXcmup1/MX4k/Jgt9e5pwf
GgsgMDJi6SLNGWncbfqFG17BI9xT+97n7tK6qBZpmCOf13T3oIavJYe92dOOl1jQkra+YfBOgzfs
5yaIt9CQ5Y0KI8/MzRPPw+EHt/rzQiKJB0br1f7e6Od4nqAQPop4+3i38MwubwkxmuY0Nm/ztjl3
YwaphEcua3x4KDEtx9peBvKkL9DSjEB/qUs53XtUb7zo+C9ZrI/9in4w95IGn1JF9B5OgMriwu1k
nHWMls9/VvVjZ4farcqRfJxkmfE6sA31T5qkZ5YwmLpj0JYMXKLucnqzZ93o2D570acVP6fgFgYX
qJYMW733XgejDn+SmAMnlYxslHAGpUA9NBEfYfM6nvyAs82o76TLMZbUbswaX9R5nxCqdYG9GGdv
ciOkaI4uVx7JYdraD1V0EvTip1PH/Ne2CRqcLw2oZPQkGdROBIS0ZX7Ln8Sa6JaXHy3/1iFSavSP
ehd3UxXD9MZoXn1nu+B+9w4iI5ct+2HnDi+tz7MlXOHYRpw0ybeZcr+5ljjGhIMJ/cpMWrmKF4gZ
A5LrA3bkwrpJG0UryncqWb09juJ4shEH3O1v1bSNGGBgV/Vxl9gR8CgyAu9FT4p83Ymz9Rx/pbWW
bhX93ZTg3CZvH+YDtHyIb3VokE7ymhSdiQHLMKhkPzXURmS3Ar9l6Tkheeqmy5uYnIlxDO9Z4lmn
G2LInbkMW0dsNxA/o0xz4LbqdWw/ZmDjAfgnb8JmHNz8OCsx6IsjRvUOLuk+oFI6hmXp4vaEAjEI
jqy96i2U2QMfYwSZJ6RcS1FdIIgkxGia1Fo5eeTsmZ2CABgvaFkI69jxJTUGPDC9WiLLiQ+vGEi5
pveo1Wle/Ey3+LPNaLfU6KXboYXe05YkA+BhFT+7CXVZN0OqIuWc6cxoeiZfVMee0PD1qXUwpviE
2GtMOnPFgH7GCDbTEDXivwLTlIYnJNqreBdbI5HGPWkwfid1RzGUY3GkacITtLrstQ4FuHPHhZ/n
RCo4XAUKYajSFkFfL+ffgF0CdKw6De/dy08hU4o5Mp2lEPbu0pU7Qt0FkvPrghdugy4om/n8DR3I
u2z9qPrd1vQBCQeaAtrWXXaydRP+dCJqM6FZOzvothLL/ygAn+g1x4kI+QT/YdrQSY1GzGXwof5s
NN5Hus2K4Lkpi3cFo2JaCnT6O5fxg6wB+PmcA3Eg5pCsaoXXixLatEzy9YA2CfJxus8NU/wjvuK6
RTgDCA/D+XRPCxuTAPwTbkM6wkv+gpDNae2JJ2hjFUrn6WLsJ/XNh0/JAAqIE1mnAxpoW/aqJYxE
T+5NpdeaqXFhi+9VPiuf6FsqHmNBUsNHXJrQwx51BFFAqYCaAxMhD3yCUTVQ+Eyterr+2mglM2ej
wikLEkY1DOO1ixYI6LS25HEQ+WLpk7NQcFocbJUiAdvlczxFGgxsthyINBQ6WC4Yd1sTSJe3wy0b
GUCvQ3L2MB9cnB4NxnkwOYO7vsDi/2pgyGUCiyxr3zpY46AeFn5iQmlSP5sKvbPoAbsRS05CiDz5
YVGa4EeYOPZNj5wBb7d4X0Ksumotb/j4sWoMwpru+TysHMwKhoSqIG+rxb8CpeAq4DgmwesFKoLx
Qxfnf8dZ6L1V2wSdU0jJkkgIfvutSjhEMCxqpGr/yixwcQT6NdDA5K0++eOs136zQlqZjselHcr4
pi0BlEg4f8X0KL9ITCFzLhoeW8Psy2IYx2h31DvCXiXIm7MvtIY5dT3CpsYGhf28PH4yEJRyc+aO
mdjWmTLcP/KNzO7YO/dLUtAUWIzNEOECcDlJl37+xakpGDb9VGAqUnScnaSow2sJ8h1pyz4HhYGj
oZmD1ssvn4gn1fU9c9wWl8YyUUMKxFM1JRNxhPfO6D7kUMZt5dyFQaTvt/DCR4Z37vt35xjnUBFS
VpduSEZvb5JeajE2YY5hVdYAJKrlCVQSFuFf2n2rgkfEHkuv8B93f6h1cbWhDHQlaGQRThqRCUn8
py3Yv6/mr7owI0lN+PGQFN3O1G91D9XsAKyww817b4uUYUR/wQzt74ZwlMmVFEWu/ui0gXsLuosV
tpI0pRoGDBbGREQIrwFJ2eG6dCU3LgCkd5AGPRRyNBNR/ajY14O/iAlbvOPjgojofGv6i2S+L9Mf
IF9UyrG4N/CPQUEtCs1mOLMg5cCpcJxmcT17Od8CdBvuH92Cnse/FLMtF04MekwWFsjWatEmFiJR
ahWnDyqnsYQZcR7Bcs+1RJcLA46hEz7F8TvZV5qZeRyc0cxylURpJhmmD2NvRKwD6Xyw6RNPCwwp
G1+zrWlgGyQp1Ovmty+7L9qZv4+UvbU4qBIObMh5xujWlaTCw9Ak8GwBcyA3jPmA4onA8NVo/Neo
yUSIbwrkBXJaG2hAAwjvME+L8e8/JrnsoLxg6ZB0yNFuXqkxR57xrDogdHttspZ2hXbSfIdc4kZv
OIonSpvNWBPQ8p8ySZIoa+B5ETrVgY/Fk4X/7nj4pDf8N6IUAOhCIb71/PzCNmOjzFkkarSEYLwV
1GV7WJj/XH0fu/GgVYpoq43Dt2KRmu7O8WMr0mHFDdtHmWeaMIjcZtU8LjIHNhndoMNA++Q+u3oA
3uiTeyLRELzMDyRVXTC1xRaYRYYkEHn9kn83Sw3U+Almn9xHBw1k5VtHRQS7cnbw6/8jjkmZT9Kj
6wZ1XEyWKbMWWnWKDf0YGlZybHWmXey6f6at1x3hzhj66rC6JNGztPM1IIPfhH4EBkfb9bhg5poz
LBiAVmBcBqxz56Xn7utEGHQ4rrGXkq8b7i2G8s2tb63LJIWc2YjB10O06sp8Js++LXYosLN+DSuD
l4GSJKbYgnqLhw3DdpRikqW5R9qzS9rdrtHYNIf7K2Y4kekpIC3o3afNhd+N5i22hIuiZa/KFgAe
g4rYo94/iO+ez1Bw+e5GmMCKZ0VMkMpF7a/91xZ469QQ2AV1qLwtyKaDEuq8sM/dINa82GzpXrgb
AXEHRndEUEII1jyv7Sch1nLIZdTlaseYltRL1e+PXZ9Q/zpAIyTsW+9RwpE4qELSwRv2f7Twqsvr
EUyD9AEAtONezsIAifQQVykJqELMOK5xqOb1tumF4Ipc3VEQOiA6b7oMAYrsOvMQ3r+E2kTrwRzS
pps/vSBI5E7vzI6dhvKIb4A80tfmPRKRWcRot4Hw+ggLhGy3NDF1s7+ptji4VNCtIcJkafqPVgpJ
S9F/lY0QDCe2+6BF7vBN7kudjxB6taMGrWlqR/DLu+q7X3SO+6QJPXesjvag7KBilsLL5TsF/My6
jcNfhYZgArD58j2Qcz18hniBYS5dPW5izUfSIwkhp0l0O2qbzsjtcjSqBd+Ye6HJm8ISf0a5Eed7
wdwF0Y2kOWhqvn1WRM2xF4gPae1Y30y/3zrX4lpaHMYe/Bf73O2zcSDGayUIldHxa4vV9M4pyXp1
CLx9rZNR6UmMQp5fbNf3+9DVx0TNQx27GiuxCMVCDbDewJ2xDgP15JldHp9RKfa/bf0b2Dd1N+uc
5vBui8b3x/DLmgVkyXhb/6n6ylQtQn+IhoqRluHMxwnKUyKMRqEUlDh6pOkruxeOX9B/cIGTPHEG
6/6GMOS7Px9ifw1BWsVGYCj8XMh2qWDNQrrKKdMKdlqT0Vmhsk2Ri9qZcydCPb/JNgNhT8iawT5L
cJVqN2Edn8PRfHeJUlgNWg1m484o6h45nYazsZLsJc6fHOLDZkNsJ/F1leM2m3u9+JZrSuC4qoUX
LZEKrpGqoXZYwO7klS9isAhoDmY5DlDcwoE5FxGdtobaEDPioaDYi69tFfpx38izTg1NWGaCWarc
QWdmN/mP6KP4ZkCqXGpqt58BGQ+egnK0eE39fYhTtVoXQODh0Wp+44YEOtGAR+jlpSYdwYnWuk/8
zd69g202HeRW+a9jh6gt2NhhaGn0BKnUNqokl9h6ZtjMY1xNBk4OCS5X3Uev0q5CU1WezsjNdvaQ
nwJzJFpC49XLlIhrU/mxRElluosjsDtTwsLMonzTh6JA5m2v4HFIOJXvx7MwR0hHcE8T2C60pubR
Z5B0xjltWgDJYTbZxXwcHTJ6srKzBIRigIh3OGMO6VWYl8en6bUwp9Klhf27au9zoakPpYf1VPUm
HT2ljsb5f/2n8AhQS6a9+8OhMHvNaVavYmaLufCWLOOOMIZcZIwfSyoq6hFmc7ybtiWPQ7aVewtj
0ZbUrByV5/FXaQQYnaTohSmpgwH7P/PpdrC/ZPUpTzIMm6zsdJPpPay6zU8RxvYYORzusvoo0v4A
zY8MGb7NiPnlyYJ/1RA7W4WyL7BoQ2oGucPLfDUFvEsmdTrHSPaUlhHzwSpD44gnGgVf47FAppKp
b6FewZGTWgOzQHfwm1c3GlVtNMhxkzoJfeqGlXf0zShbXMiwBhdEfiHT+9GT1Q/xRSXtSM5v77j9
11LMWZCa9ImJbTg168ryiiapuK30EhgP5KWyVHBT1/zHKGe3jkXmS0J60qsciDK4ilRyMHF5ep72
BDOqEcWYQj2I8iUQoZekI4mrs3eKhZAGYTjCYhkCH6jDEla/Fy0a+hKhWUnspNVVgmVimuPCZgx0
2wj6rWWEIr0C9UwCtEgkPsQufEQDUPrM+b5k64ltOhQDqJjkQ/yKL26aNdyCwfcFETkiv5Xpftfo
5WPViJ9E8aJe1qE+SuAIAbxXkrwnxeZFAfC+s25wxSPAQ8t7gyAMjliaHPncAgnfueL1yE9IBBUy
LDl5Lz3jptAQTDsPq4xhopu1OXH11JazqCNGHMkr29iCVwsARbS3ixuqPmg3tz3084z4tppQf8zW
te6Ia7rKfFugK+UAOgGOAfGrBchwypQGG2wrcK4GhX0zOU6RtsSulF3xMppGIwJ1GqnEBg1OBsgD
bqBXmwXUyhsKj04Oo3nffOEtU9snPi9knfE4J2qX6RM56K2TFA48LVK+7gH1YkTKdcJA08pzHJL7
Y9UpktEuVdyUnW/qWmnuVLwfAn51sHzTmHuYD6SqC7iY8CBZRNvVsF6VuPVQ9v1YjqrFbRSQMJeP
dfCpA7Uj0/KV+0BxFmhVL5IL8nYUjzJWZLoqrgmRhvrEhnaxDXO2SybjtEdnLdLqq8n7ppj091nT
2tfnuZuDdqarAN0ZVOzoBrYASmKojji7lAoZ0lQtCuLwWht0bbCCTV5kDqyA9OgFXlZ4X4TmOqPY
hAAB6J/ikbPZqXy9mcF7yP/jMNpbOHkCAfASqK+uUOMMFL9SEpvn6HuyhLY4WJjCPFOltnNwJAJc
65PkzIOzYYQ4ol9ZVkuhNAdyWOGz2yIcdZ032TF9FLb9n+kstojzIQwcuW+bg4a1/kRU15hufBfG
bockyyXtiT4IWSWgB5uuPoglUVx9XIIzc0cQ23frBTglwG4BxdXNXtHJewT0wdMbs3eBaPQKf6hQ
vcEkO3r80tAfDQ7sPhPDL246A3T/kx70IZKEGK5VKbQOw1QA4czoaGe5Tz/7dpbfFjWw+xyYbJjX
KL8EUvddTEUxpLEsLd+TL6ecP/1WdVgtOLzIbIhv0HE6bIuV+z8onPfR255lqbNmWVDTzo1/Lru1
rDd0lHUt5vVjM75NG7m9LFEIq6AslSDb7Qo3v3jezVanaqss1m70uYtxksG3osYbEly+tTW9MgTg
sp/SGJxdCfedk+PYekxnkNOrNXbcWbYalSsEKsdehbhYY3QGi6gTWw7kA4ys97ufsmznRica9/JB
dyX+sHOmkwamPNXiMEjHrXtY9vqy9+khQJ8NUWaK0mOaWxMHhrKMFg5ZWHyhlAWk9t3/2fQWb/8e
qC7dnUk8UTX+GdpoDwAdoWlVt67kAz1Gld8IXRRxt+uNXgmhf308UKaXMpH1gZJi5yd0ttBJQAqV
q5oB+ljQr103/cpKRs8OSu7aFr0T7ySLm4Y+kYfjn6jMRpNfwk7+cJC+87CFtI7VEXdYZm6gC4J/
lIIAi+HMxs5dsEaYiIVj7s2moU2N2PVsCQDc/yaqQJs2qEgHVdk3vB+jlTxIPCTr4/cBk74pvdcm
d+p+ho9MZzHKV2wjdZQ1UtTPCqW4hGnxJXEYrPe05W8fiFOjJFNVq3JmPQV5trF35JDErhbQEoD6
BekuVNLbB5TPnr9HpDJiG3S7sTglxk9EqRW2rNGSl20gwwRclL+fwriG47rdwlNMVfOFDpTReYs5
cOkte7MxpnGlXxnDDsVmMflR+P6duc3pKUB6vuypiWCZ06Y98eOJTXZv/OgVZNC3m+Q0eMOMMi7m
CQjp9r87dHc/P9RVO7AR42sXQnub/t2nIm2+ADpw1ZPo1oIzZdLF4BDzTUeEm/ZHdSdyDEs7lQTE
v3lPRkrYBxKgmHFRivmoIE3YN7ROTCjMZwum4MMR3EvYL2mGQTo4WQa6nxGNO8lcIVVznFMJOqOn
g8zt+9Q+NvmEej2IS9KRSRa46DNpDyovXdvViQTD4WwMrtJfA/18I+/878Z63O6bvnKjtACpAwzj
QCc9RoaBAVxx0Rzdf1AnZo6m14SRiRyZ4yeh35CYupYUseL4heoXvjvJKiuYuHKW/Rv7N7uExgZZ
CYz/5RUmbWotJSmp+R+Ft/PtaqB155s1Se4xgEjHLitTGnv4YYkUB15hkG8DON5RWBJTcwFVyzhi
4QdNTP8TReJbNAqdddDk4RL7KSCOSOcPVJmZ+LQP+wAd+KKamqpN61uUUq6zfDHg5y1/sAVxSYS1
HV3s6ccPRfxMmY8erWfW3hSQy3GHB1L8A3wrVBzkPJuy2sAiBs98ANBkZov7XAO1G42LBcHgp1s8
B6AtGDfBo5PMEmXf6BnHC4KiGvwXS6KDmY3oNY9qzXA3x2v2tuSoMurvaRhQh3YMDkQglh0Sz5xb
O88HKohhHf98yHczhejQ0fKZPUK24F3X1UDyGXdZdvuipSBsnzAkeQ8ngswCmbv9ixW9vQZDh5lx
k0ONLYWTy0Ri7nuf78EfVKt8mT2IP2k/84cUKw6vSo2TMUdPbpTN4xDuhmSKCKEbcaDvY3x7EFhU
mFNSYMBtcdfVvZukLjBiKgfq6C3MGmcpjI+ldZtU/yD4AceQZZuRK226KK+8sxM+9MlIiwmdmVFE
sOC3j7q2Viv3My9lLYvEZ3cubK7A/JFoJ4IFoenSYHbHay0vXqFQjIka37yrApHEA5LMnMNeCTY5
0E2G/bKS3y+lxIesgc+hl3baDe3gqOlC06ezlxsTN/7oPcm6KnwRtdflMxOBCXliL6I0eCsCKXN2
AEzLRjW2eRk28tuT5uvArTGGE7M9J37jqyGsvqWGySC0euysoPSSv7L7TZXgWdTnzdoB930raIwD
cQuNhUgqggWlq7mHTMFamV5Zn7qM0LIB3ae6R4N/Kcw8trLsbjl14/MxUv7ikqTVI7pigCFm7u5c
OToXiV7GpbuloucdFXKKTH346v88TzkWHgGJQcZIZUijVrz8XptuBIKq/YMHYju8POeApP69zlOH
Wz0EiqiBq9apr8EXOE0AXVVg2qZw//cA3o84qbcpvKZF8LP+UD+eP+2JQd3xPpZJdzINilzbDt1j
3BHwjZoHbSbIjsmTsqNcKDpQ73ZEA2N/Lkh6UXiR3WZsSHQsHHiC2g2EpXnCVQuSyhP8shXntu3O
S/n814oFuD+8610aCi4zYB4j/l3lA6h161m1ecDxtzGMF8bRQWHmoZolqwv6zHEKlpXgaDPPPR1A
GwzGE3Uy++Q28t0tab4Z+B90XefER1fL0gjf5ZdVfHGsNq5dmzjjPJVaHVXdvff+Ltd3VtIxNgtD
/R57Sc9WFqr+WJ8ylNSWVeo5wxLjGQtbC742f6u9CxoyBVQlJ8UVX9iLJqknMMgdFNMVs5V/Uc9p
nIICLOdpCYIXWI0ByvhYeKdgakuBRIlfjftEw50no0cLcKS6jYWRNh7SqnFosNbaQ67kY1RtXgpA
f139JDpppRnK5Kg8hAOLqrhFDPFzikkH9DRXImA4ci9sSn3hperba4QQYNHHd4G8P9yOmd/DOJCf
H2OKf0YNUGt3BCl7XEhlmZVEwiRk9v/nWN8kj6vn3wVBd6l9H8xeqEJH3BKQbvJ2lVJk1ZU/apkI
WjksVWSfg/VReo+OuKJQbjU/KhWbnDZz9j2o2VHhSvLtapVNKEzs6oUnGgxxGEpcHMUWyn9ngDrg
K3ioX46B5iPHBODDwZ+B+pt06vSizDctFcCsGVA+Fo3v9pObCnJNimbkEPsNS8j9slVmaNFh9PVE
MpDmEmwQ9FORIyCstuTwzHBrjhiUzAY1iZ1b3YkvDBsp1TDPM70Kqbu7b5x655NSAabWMCd4z234
xvjzIX/HeI+TubwhLiL7YB4red70kJRaKcHOf0pwZqgKynNrrlzEvpjIskrAE247aDmTkvCBaNM4
k1MtSkBmEBRhjA7eQLkxZ0w6oEM20uFcP8yucdBmXTZuJp1+HADOfzZfECz+IykRoCM612tLPn80
ukry/yPWG7A9M2b0Z0uBnXVuK2BdpV2RcEe69Lx8ZtAy45KPYIVKmypK7z2YaTybANdwRQ4UxgP0
gfZSJAjTJuSmX2HKmWUbsFgrMXd4/xhnGmvh5Vspupf8m4a/Rb5avdQn/27dh+seCWGl5HH6WcDU
N9kK0jVCrbdH7iYKoRPCBUxPvO+xnVh4YISo4YaoKByKHfG29n6HF0/4Wu6ezuhvmmYpwitR3Q1O
xQqYfUlqXG+RIDgifB+2jpr8YhINvHzx1sjR+3QxzYPwXWeNu5Le7D8Yb50UtJoChvJ5mCo1F4Qn
tblqH7aLrh/xv/PwTeEdfuMSuuYcazIibFCO2AxwAy83w24StV0xXt8DuVSonnivpoVoZANE1iY5
BtPhOWywhfdIn9wMbFTx9u/DIa8sgcl4Zra/xOdkIuxWZ5bKzFURC5U08SUwm7pLiD9N2DNBKxF9
AlAyMyF8CkuoNrM0UrY8V6dbnR4nFj7pVvWfPuhc7vT6c58xSaI0ZT+isrBY8vOrWwMO0scWEAPJ
LvZxl+q/eTL3nYz0gOzqCHP/HBFup/1PHfTeespR/fLTWWIXUuzzGitgNA6bIqNC6kjlJC1/9Atd
C9MzeIdKwFVc3mvkJsyF8n8yL4xKY78L+G+f2oxWRwxH6c2mpdqQIvp2RCCvwidFZdFbtSaC9iry
7dKj4E6rZexAKYC/WoQ2B/7u4PDbgrB1rlRJCOm+O9SdQGUgRjWQWLhN0fRD9baTtLCglvs4etD4
XFAVlNcMSx85Hsby6ogB5tNPmqYOC2MPghi+Ahb4CIAwITP/d93EhfMjFxKtgaHNgKG7PA7yorcL
J7nXMpBE4EHa6GL8UP4h4Y21+yb78XXdaTguZrmmcWxKTtKtHfIoxJ48xzZdAJ06pnwP8yxALkFA
mHjV+bR0m/WyY+xJPsFg+gWHh+Im3YJ3gvSHuJP2t9flEuiWwrwU0D+OTxkDq6o8MD8+nYr++G9d
d8nHfFC363J1Yci0cUzJoXJKfDxRIT2pc4C7mr00zndlIEAISVSaOq59IRggWf1te7jCHumQAvMr
T7rMEZLxmtW6TktfjyUZl5tYp9d1t6AerEUSaAvNo/C2P8NP7j4XcmqZZ0oB3WBj6rpKmiziDhK+
Urq/PvoxJo+9imTj8hWtwvPvydk9YrkceFUFbPdn0VelmUoln8/oeMZ+Uv7R+6hxl0dPspAp2mLx
4PXWurnk/9DK/qIoIX2buPgnooH/n2N+7Dft224rfkZuD8rlzI+rWdmlxrTN+IUZzVvQf4ZdvlC9
DI0qJB4JwvfhLTN7jq74hF7sAcWe1exGUIfV8nrTp5G32hzRmw6nLtvxGwbnzO9sVPqh+ZOIL/Au
FcikrlxiCPBE+qnKigDVcGqiDpuecivIj1FrEvgdiG0pvzbtX1qP7u9qHEnGqrsIqTuBdIr8jFuc
z2LDvRBty+biIlc6U/iyLQrYUNNt6rbwb6OKfd9i0QVN0WibB7akbuVRQd58W2Bh0ZY+gWC7V5r4
4v/smg93bRheepPmofV+Y7G8ZURh4rzIPJqJfT2o3qGQSuN1DTrOto4FF0hdpxN3QAkI4pqLhLFD
+oQXjjWnM3NSg4Yh4XkcniPSPhZVnQ51XVy6R1b2qW2a2TebJkU2KsQFID7AiXLIQkvMpHX/MYqz
cpNhuHECPysqNuNxvrygFW5KEfWf4anuslqBfawu7QdHjuE8QPa3HMQujUL+lBX88z9mGV/ZxrTR
7FpW1rpErpn+pLz+hAN/d1gew0RgPS3qvNay0N6VkupWeNsHwnx86/KiTfPBrVF0Yjim0ooktX7n
BHIbRWMx0YzcrJAZHMPFhn1N6LjzjantOdlBXrO1hc4CmvsKPdV6H0x0OtYGz9R17uY0BBFKS9Sh
JAWDK23PXhMbciCYWi3cIx4pALqoeDdgGjdV/3U+8KtSpsPlo63GaviTOqqjSS0dbItX1xTl6HU5
VlkG6C3q2g0kBsRpNt+a+9tjec1w7iJavTLzc+/3ASHRMVkgxFZQtuwDFv2vTjKiX+GW0h1AxMqp
lp6INBzY3h/ymqf5VeLJugT69ncH6VuaZpkagcaZjx4fZU3VEJJddsrKZyTV8VyhqRYVSzsiyY7k
p964xRcypVqFEyIyQLi7hBdp++63mH2AlFeAY2w1RtA73AY4T073VxKYYgVIr959BN0kUtgLenK5
rnzkGGHCTaA9j2kix5JjW4rh8O/DM3kDtsM3GJ52TUO/q2AFUqoPDDZZqn5+Ls07+Gwa5XTpR/Zx
cq5IFeePwuzNyzJFD5pk23s9WUVmDny9NxXPj5pegUEBTj1p5vKcFNVBqzeLM7TN+x0P+wQ3PWwc
+7ptCl/7lAxhxtgdkaUbzF9mhS8d3aAPBUdyT/w3NsheuPTpGauKrhzDM2UJY2BTzlG9lIpa3ZcQ
S+sNaZ+NaDDeMnz3xUrsk1Dj53q+Ip+gR5I0GsEJdpcpmH/gTU9uQwV44GwMPFrCsrTnJu1F8yzO
MXvxxRPpadESIKQOT4UlKSGeNY+k4G71BAQMjmnoHoDHSAUGQFcg3n91XSoBEncw3+VaNFUYN/Nq
Fwd0jypSszsOqgYxNCC5RVi1Du6yO47blYeYt2AS/6xE8ErTyALepN07x4BVZiR6Z/xoPyUcKDxq
XfCEWaQdb7tBtY46XyZPmCxBmGbzl6S4AygfER4SfCHCP/xpx67CqctSWZ3gw1P/kBKjJi0rsU/A
JJ3RQO/LhVoT1o72MKsv9WyOoZcin+JKwu9U28wW/gogxPmHzCG0Du4C0Rx9XaAJfll2fVPZVCik
m0d0h1VbQsOO1ue8LyXa98w1j7M01HtqnTRPJvSbOAqCLpHLxntQctd7SpVAOvnFetYTj5SvWAmX
bhL9+Cx9abFbBmDLPnzglCH2jgb2mO1KMVw5z1+VsrwGMl7RwHmYKlu1RpyjQQxJZtYUjFH0DuVC
9ItdAAqNq271R27ZjiCIkv9V7KA7i5JgA8wL58UAKyR7j9up5WPDpeYV1+tdyrhFSUtZK6wJqqHp
e0jL1ZLGeo4VdGjWVQx8zatxs/fSjax2A/ACoUHI6/yf85vdJ2uZXcaxgaTkQt7gHLOBEFXswgOv
WVfP0wMotYVsIQUw8QqAcQuiEXmpkKwT3SMWYmSArmYaM7B5PW52H/40+GfcCCiKjgwfhxGusuov
lj8EgKbWtWIqBwPlzpFftNjJgNC4IEpNt758c2BrwACPAYhzTZs4ISQ0z4h0iZvO85/+OvkjKGad
vLTz44cvjlrl+wL16hT/EBl9Ex5M7I6OYJtnbWbosT+gB1/fwCdJLVIsfmHX1gVo8dQ4F2uyRKuC
jPjJZK78L82gXcWg6Lacl8wk1IQJm6UTTM0SUt3zjPXpLr9+GjyIIa8QKmvVMNnWPPzYchvA3uLi
4AcS80wVpiRdEwfFHgTpuDA6UfIhePlm3ZE6ouYkgxv42Cc5Dyi10YM6qEtUWj0lO9YEoIg5IhnX
GFVQnTQojKNuUkLvXLvOkv6SV+cqoF3lS4iH0u49iBdL4pzvDhMocTkKPLLznzbuCqJZQYhyuO/d
XBHBwjEvnF2l2JQsotdgKZYqNOEm6W9QrMdZD01EDcr0H/fPeDXfmNrCtJ7MykaJVjuPgA8yzaAM
PWoEYzToMhMISh85FH6qN3TGfsfaBPckOJcBNSPUvGShIxWFLp/rCDQS7Y0IsHNgTLy0mat3cNSz
/5pnK43G9BB087On3GJf0RWln9FRkI1yum9jQiMIbn3v5H8OOQvYw1xvdbd14yLCbkofc7cB7w7F
6r+k+sLFeBIx+FTODHEaz2zystpGGWFDQBhKQizjpjciVwqcs6HcBxRkSulYphWJcFa50nYiR+Q6
Eqxkyqn8M5ueBPt4rsrUU5kcDLljJzIrHC+LCQO7sSJJP/EX3HWGIg2UATGdmTxDVjjqE9poJFg1
l3f7DtUy9rNbJWRcrP88+CFzOhdhBn26YqpkA86kDDuxNI/AmWruHVNy83pwtjfbmQAXgfTdJAcg
7HdUIKfSgQhP4GxSOjthUVAENhhdVVnSRHmZd6pc0FxRkNUBIz4jKd23k2L8VEHs8NGU+36CWdag
jvKnj5XP7uVwpY7/y6mQQFUMZsGoYBR0Uor6w3t3wURtQYDngC1FfVBZeTbsFeb0z5IF7b3oBxQM
qD1ykBglgDGEutQe7cdFziw70U1KELLKv0u2gQYVRhJK9WDYG9R67/DVf2TcNbEr3iYdoSjcjTKL
pnvImAKui8qYu5WgmJwCcXaW0My89KiIaKtC5yKo780KSwyAEdsFsAgA6sJcYxmYdsIxSxeqzmy8
WtCfC3a0Zzeug12kz4+EI01+ZppLQuQ7bqQZjte+N3Wnqao4TdX6KE+VkoXiltTD3tLHDoEEdHqz
KcJaRlEfd7MNQh7ox7j5vGosktKRzUUaKU/WUlKBQ1VTou7pZKGm1kPIsOOTWrWsB99x5FAUgr5S
C5sPWIZKM1vIiiu3RQtreXLkYKkfdczb6HIJHjbfXSuoHqn6PBPmLEaGGDM/IEk42SH8tIuKaYt2
KJj2L+nmKpR50py+xXtM/sxb1QkIVr9KdtLqlcOw1TwxDiuqgFeuPQZDG/T9MrdhNtXmoJTJOmMJ
FIe0Urr1A9V33f+2yJ71jana7L8xGLmGek6qIOLjPnEeRq3aBYm3hEGQvvH4QlJf0vzRVqtYxMzM
LYp35VylM571AUIBCYKoby4Zbi7c1DdY/SrIf35hLgnOqWEBYeZNu93H6QmPtZUQPvLk3+1R8oqH
pMGkSimDjaYZwb+buJYcjC61Sdb72JMyw4pKlhv0sFEJmhkMicID2FQNaH18N5x3Gzv8fUah3nGo
7EqPtnHQQwQVt42oX3dQOqGWik8oIRpQHWjeTUTy1PscYucqPCEXTELBl6Q5UFml4QDi49t6mlJg
SChlhBzlX/9F3tL3eEZGS/w4yEmU96Zm4qJK9mNH3gI5fnwuH+yzWOrUM+EFsTReVhFhfCSq5TiB
ZdET5HWMOE8qRsALApxxoZ2z7PGloCAn9lSqkAmm2PNtRaZPicaElHeuFrsbdxr3Y5p+sUzcJOUf
uJ1bi7bVfOCg4Mg2YDEOvnGgN8y0zgWkCrgp81qUveTloBgx5+UJQgTRBY7vVQNDxLQ5CO9ue4Qv
ZvpbR1jBLjd5RIfkBIDRoPfwEPE38Qx1ErPJ4hSKQBhgODOpr8cQCIWh/PTY1PvecRWOMFSSFO0a
ndnALeKVpLTG+3qjhtGfVAkU5+Bnsk2RhIQEAdXdHxQcMXaadVRhPkjP4a8ensyQLzzD0ecgNRhd
QjrlvMyiOygsCjBROddb4y+1krtRAcCwSw2CyR4POy0UfCXpK+FRVvbyv3AbFSRKsyg/M981O60/
1MafN0FcaX7QUt/o48Tu/EyXTDSIqauc0Bh18hTyerEPW78cY60ww0pE+d3ho4qtrD+KSMO9Li5A
XQf2k++yhmWbs80Ec0Zd2I3W4AvpXtv9/hcyAzi1fnw7TXmjhaUdnvLQr7ozb2E8NEUnTvnEkt1j
ejWpZ10dvdayrXVAUWT5kTp0mj23V9ASOrt68ThzBt+53YuqkyliH2SXZROBb5vIS5okNgsHshqw
wZWA8Kq9apNblMyf+Zc2S/ZCwARMobnXCZj3X3zIenIe8XoakWj7oGuGaEmsXU5FSjcrgYHz2RKl
qeeYuH05cyHyUJwHRUCADmxzzT14jEtNOX3g7Fyx+kqdN9qMaJs8DzUa7KqX0V7XHqj+v4fGGxhW
fJBf4RJFjiPtIWqDcqktgkzqeSCY5plBuUOsBBqgojCREgxoF6rFG9yCFmsM8TmYIuCVs0fQIvMn
6vQKaVTohsAN3mKDfcnUjJ/yBd5khqbIa4DWJAKkSUerSNktk4uicni5AUUxFXvPbsZV+K+pAEW1
GB87M+DJttZtEtVdhtfeSh2vB8elh3FmQw/4qU9lK3oCmDhtdIJGg+pGRxvy4Z7BSKgWf4+9lDli
SQHiT2ywLQNtY+e3+QUfKMCzb4zt/ZdLYUiw7P7gwiSfJGZzMDZGl99GBdRpKwoq5vV0v2PBpaDj
mZxZgTrkmoXwaYT0kps5/1T8mSMM2ZvZQv9hipsjo+yC1jPpAw4Qx2ezIpGgX1AM5WMzSr8+uVnX
7xaTkpudkWhO0EuX00BKw95Oqg5RfGDrw8cg4h3FnUad/mZF1MZaU/Wpn37o3z0a10OQS8d0mxwW
hKZvE99F8wcPSR9FlMTNPMsS+cWI/bmiTAAzr+173WMuV3WLVo3MCbb6H9bgesYddGwYvIDsv4uY
R70ADjDfC3TSbub+vkCi8+2KLuFOMf2lIROaJJ5QabZDkjumOtT5rFCBq+s3FHxaeBlmxwNDacCY
OrXYC8jiGJHpSik401pOZoWu6aSkvha6SX0Ng+7ZlqrcJOufeIGwSupJ/MgPaEtabPsmqwB5ZwUL
QCFunQ4wn1Vnr46CFwWIZZFWOE+2fed+mFX5BXJ8/MR2gFGswymadq9qvU6aT5Lq20Ps+NY6uDLR
BHAeFtZaCBQDlKu/C2OOA0io+vc/etdd1zjqUUWN0I+b8bbSW1o4HC3+763Xoo/kHUKouqdOJnKG
4G/D0KB4fpUJVcYmUs5loDD8NC2Ky3lipCfd5ce61wggijzRXOndJBNz7hyh/tBzJvsSDsCYTWYC
jTX7sSZ51RpWRqxX51zo5E8hDMdAgxRPEm+1aqw1NI8H3i/rCWaYo1hc5UWcVc1DeWvjGzkWrAcc
8YVFUXHd0OtGZ0dhLGNOG07AP3kqKNCFJALFYYkdJygVoL6mPU9in8fKXl8EU8PM29kajMKl1eOY
L+TaI+Yrk9fyQYA5GsAnrF/l09s63n1j/v6SbvNJpgJBTmBhFGy/m4K63iIU1imGQjRAHgKOhlUT
u/r/lk8ZEKtwrkUHswKluNTIT9IKkbEsNbNKtpGtvF+Qs+Dj8OSIVh46zmjOwSi3gQi7bbby/V5r
o9n4qVGxfXU1Ut8NGa6NhatobcUZYFqna3uDef+4NKA+YxV5IkOwD0NsJFcxMw17FozUlqSaWmcY
FcSHgVZldolKTHuE1VBjRmFfgokHtKmM7lXhFA3wq/C0eQy5ZmLWSlWnRWahlmszfg+FM0+Ul20n
9jJ/zdVumn+yNHf6khCVOM0zL/hdQQ4470fZe0h3ybS5Ga6xOFJQKt+qzvtJOk+kmDqcNplBSU+w
0EpvLkiswtiVBB1qQp5xTEEcUTnUA8ulIbf26e1SoUmN16IbmSQeWa/g0JWBz+zf01nLhS8Td/ek
VimDl+snntt/NnK/jLL684yu+pC3KxDXy2B+F8yimLaR9fC2nt2gxXZABLDSKlby88lu6rzhBymQ
z3C3unW4I5ZdMzmtdV9I9+2XXakggrqjMeuQ3CbcLjpZfhLRzEEoaKkx80mJtyJwg4KFdA/5bP1w
b/zBH2A4bUQCWN1s4y1243bXa1if2hW4+nZc1F7BWntiS7scAZPzvr9nAf5T/JdlisRgMCbb4h7g
17m6dH+VpzEkclszWeT0PxvuTzrihFTD+spsL72vGYFwQzwu2kJb8JgGqpa1himh9tCne97BA5LZ
qjXNC9oSHgqnWWTv2gJR4JtkjDchQ5f1oPbe1iuQ0m8SeA3j9vDpdey0IfX95pWCQnKFCpdNfJMs
VVxmpWL1QYZFKt/WT7ryARoRz23dWI0sWUYhhYsC+RXmT9OIwb3JQkHW/+k9MGl2iHlOas/gDe5h
d5MD30dmvDTfpUyZ6pGtjmj6elLMbu1UXgEMVyvNaLXBtTE9q9fpVeCGXfoLzUUfC6sM8ywCEj5n
ffnEN+4TF0gOgRxlsUNCl7wg2yfc4Z6IUfwnDhqM195MVPvORc9xHLEHTJOSzVkaPQx4bgh4V7YZ
nEgUi0Sh3nd1LmQs+M9Wg/bWXYb+LsYNZHTNkeNf8tU5Si9zAtn4BjVHHZuj/C1J6g5zskGBGFEh
eEN867Zng01ibkASC4HrJTmE5pd58aLO8wCT2Dnl6BeUyXXgaClNJRfi8g+BcS+ecG3KfBmYaUbu
cerBrtDOFcTa1Dbp5AzJxH/VikwWMy1wdYN2Eo4T+zyGdYdtXueaF1wgt+Q7nSzu0PP4w9KKX5jq
TgFn8+Ejmo4kuatNiVYMffStIgT7tNqo7rL9jwivBmLJcg+6w/cKUKYAkWlWCfMZ4X7/3CqKK+Vr
PFlv75ov8ft9NSGAO1UhsDwnfK4zXgbHx+fth8IlPFuZjQKtII/aVGZ1EArgyJOP4Mu2uoglpslq
jlWVKwJTF6o6uIg5FyODSUmDULXe7WCIp3/4E9oRR4Y0NyTLjf+u8hcVLfH1DPs6RLmdDbzWdmJn
HY5dovgQfc/L64C+ZVxJ89kgVKCCqJasGuvpRIqDyy9Uj9icC8ime4n3nUumUgygq+02oQ8exEu1
jQlSuo56JGx8TW2/ymzlvIN50VlTaotwgBx3lnRjp04L6KMlcJw7EYOZfOu1T+xdutW65dW/wlOM
XQca0ouRE9RCaa4H//ZbCFjf/FY/V/nS35uWGmixFX+XXH7Sf6GCRhc7GpWGEQnbgiiPTd+tt1AQ
UHQ2GPK9+PclpHOWM2K9wKRJtC6pOAwC3CiII76fq2/cLuv8KqNem+pxFkVsbN68OdV0hEzG2Wkv
uBOGZlxq0VPvjCmhvDXndBjE9Q+0NXJaN6EOEjOMvSzoPbBsq100l4mahJr8QZoTvbT/yVsReXA7
RrXb/SNn1GTPcXsQYI0atlMA9gfSBH0uHPy5Ag1Fi1RcRLxigTnWvuF7AIFTe7O9N3r8FYb2pAJ6
6TRazedsDc+bsxU4zKx2Er4YqVJLMkQxlLCF0dNA0aL+cajV3Ox3jCyEB73c2NMsJkHPpDUz5e7s
wyov306AVzBiku9zSE8CLQgXFVG9hnzUJ0t+YcU6osg7KadJb8Qs9imvF6zRyBljVyE2RGWxNsEP
kJIlsYtv23PYqsev1xP0T3MI8TaJTgoxaPfsZqMk0mti4Eo2DJua38iBDSRTjJgo83fooMMOv3br
WcD44KtEmCv+n8V+o71+Iwgn60KKKuVnLPTi4jjDVR8bG+iKhUAE17sWW2ElQOiWCv56LDudvFCd
ehhk/IzgekThe+iCJb0iQixJPJzWtvp1pTRrK2hCHpiHTNpdGnP1+a5vxT0l4tCzr0Hbq4SfVYN5
44yBUnf4dJjaq4Ll2jCuAUSCeA1D/fzlKng6A7HnzZJqKjZqdPndadXd7l811tETsYQYyMxHn6Az
BOsDWyGavcAiEXbld0n47Ipdq+N9mqY61Tr+GDJBJ6viZd48gO3M41lsOiqvNJiL1ocKmoglGsQE
TnFiCh2A40cMAIxZGVPdAqS487iPB8fMeBeSer01bI2lP81AulRLpsCCb0sDo3BIFn9DGhEL7Ly7
lwmuh4WTziK30FIxrNrSM4i9GW3LShNE78GignoA5QSHMuRec+1b3ycqwdIuoBVkiBDm5xemfm9+
kEcGq+hIsJ5hCLqXwyBp5E9YyVZ0YZy9VMYtLnD4NzJpdYYWL7DSzsaBX8Gjd/0RkmwB0dCKRA/5
/XQVzKWRwQWA6rlQBezVvtkRsbfBK7qtF3tN06cA3+CfBTIGzSYtgWwWVSeMYddsTKFXLenWcH0I
5DYe7pXbUxKsWdHYwV59q1aRIStFXFcTLHBz4sLKglfgOsAp7o43nskeLwXVHny6FN3MObG1G7Ae
o3XmWgzkpITO1Lo+TZ3b9xp69x8OeM4/CmhCzkd3xv6OVgbidYjIvpg5etzKhe7DqHV/nIS4Npg3
xVT8PdRzs3CzqqBgRCpWBBlfCWDV6yLzGjda3zygFrrz3ypBHeQ2zKC5Gm9qpS+0LbYiqfmt8vxT
UND3PXXgLuAEWxu/1f1aaW/36S3lbyv666dEwmoiTAcNJt/Y+tH87FYx/8hYwPlCm6XJI+ttqs2U
EJ5wvLx17AsP06P7OFRjrtLiC0wss8qfRZynquUH7VjO2e8UpYbsWHcw0+zoq/EY8TbrbQw/vphA
4fKWWIpXh+H23tDInvv/8EVkfjpKT6/FWhqo1hKvUQywfvnHzH7Kz1PbEKQJMFM88sCl4RSQjwaZ
7s6lAIfNkd1AjD+OibCCkWviaoB8cy1wzDj/6SSMUzKybFG/HrPGMFGgtkNsAWfC49yciVWggBF4
N/yX/782jTgWm4VLWHbHEq46vkx9AVZDGRs+YTxn+2k6BWPzupiU2K5ztWZ5m9G9MJmNqbnFXVnN
EiZ7sM1Y8JgoS/yAVonAhBY1FSKuVDsfxagJwZW24i91lnAI/A8mHm9fMMPd+aIIc6hZEI4Ofa9m
4n62ZkNeQrn/u9bOzQFllbm+x9uK7exVAapvnPB3/pqhWumi59xubHakh2vz3pqmtAJOCPn9s1zY
aiBddbZeV6+lp+ZaOy5bqhR3w/973XS+mANTZ/AJvrPukBR09RFKVNLvtq60FHUsqYQumQMyBRSq
KsNf9Oq0LTdHlY8k1P6o0aQd9PK7X8ku/Q1elEXkxPFIw9oqJkqqybHys0KS3kfJKGFxocFmsL5Y
R9y5WVx2oJ6W901+rlPNg81Ns69OpE5KHdujC59RzOtjdl10M+0lGWwfdKJIunvDCqPgyQijEWxE
pNkyqIbINIRdqEwTkhcqi8QDwr1Klu5z0xHVcJaS+eVEadqB5U4fV6vLOUHe5clx8InDZDT9laEG
C3zV4Xm2DrKgV2ZPbgO/JijyV+aa0Anzet/VyQ5l/z7VMSAMlNpphStcikHVF8XWzFyhoV25TKk3
krW5da5NhIbSqxZVk3VFkEp5qPvAjM8HBnGRleOsV40zAVgJIOMlLFRDEHgt7eHvU2Ru7ZzMepjY
5soz+gcaJjYA2MQLNIGu6soFO9VdYHqFeModpKoVrsKsPg+MeCajJFNymye/R1aIiEdXvG4sfulf
gsyseoLH93db3ZUBO8AzkHOKjLr/q2y/urxkXqL75KHtRa7MQzEs/21m59revGwQYtNdlXGT/exw
qNnuOB9y9iYnircIZgJyPzQII4nll3qp7DcEfz36kSx2P4nslvWxPlK72IchmfsYV+jPV7EkES0J
lYzEjeP4yjScdwBvvMK220k/qIVo+fI4XtQgd704zPc3TbiicRqwOamO+2FaVxXcwk/WJDiwZAlF
GAhlc/njHIxD6zMMEnG4Iowb19j+5UE86nw09uyQgkdWyvmRZbVgNjzfoygBWst/RQBbR+qFcFt2
sB8uQG6vOoWLlUjn2EI742NJuI6CrDD1lPnf2LYMBTAtGvHPAZfq0YUIGOYUWqV0sAvtkRspQol4
HczM7hmc2nJguPOZqpI+EBqawjz9DOSH9Untxbknt8v4KYD9t3vEZKiBbX4RK99FLG4L/7ZousUb
qUQsjJeJs5Dm6DNKxbEPH5RZTSzeAcgThTZGNFXlPcZyd6jN7TGwMismQ2f5m5UUkAVSE/DqOwtx
s2AYzeKMfprFTQ487lTH9CVT0z4kEWc2f0du+Nmg8gh9EVBh9Sg4fJ30gOiDen8PbqMz102xLN6u
hhJf0hSGHtL7ETaE3ONVX1BrCcPNJWhvQ0uSSgndXAlcHsVl5+MpewF8rMB1s+wJkIeUx9uBaMhE
h9xThTG7oMRFaGMitLnFHf8JB+DmXK3VFVr2gI/60eOELKcS/DshJB83xmR6qiIjN8rPMUlozXY+
k3iQTBvCfjlNNwsfBuJymg94tJOcua9XYq7Dj+3kJYvPdWAC/+D//+0azTNqjM38lojEu+0DL83R
nefymF1/9nvLbnoNOu0fNghkEhvOUWbvIho5DMeSXwmumiqeLDK+v+OATfxfIVOkEOBJfzJbbQJp
TYhEY2S1VaKPNyg2ZhX+dDkpn2SpZvbygTmm/Z6z6Xf9sPpCqR2tWWzPpwymPVp/bDYTyY20nSex
ywJj0nYbzTzb7YVFHJMNruduJGsXIrN3WtSZbJ0+xaXC02NkDKALxI2XNpKH6H2nXibkCKdp09mz
7cUk6C31sh/SOHbr9EuKzTa9IVGihXKA6Q5TpTz1kZw0grFNnSdNvR+tmkIR/bkfFbyP5BdJmwrV
VPdXBCEg50GY7LqPlZzmgAeHRXzzetx8g8ujTGkRQJnzFE9MUlGC/Zc5lmkfRo+3C0cOen7riioB
RbIzgf9nMWExAgYXE9/XganN6Tf2zoEqn/6xlbiPwm3WTspDg0N1E6UVneJka9MyoSFPSy3iibmA
lheLCAgHAPT6KI5EIcG/HPQUUEE6t8WhJrY/AyuCYF4iG9O3CSlnr5GQTieyWlTmxMP1fqnP6mC8
RXahjrEIYFp55cEH1oNUaKZB1AeCgyRksT3a5Quov8n4qNlPZ8MTQZCf0a9KFXS/JKMY8LMbP3VW
uurn77m4aEOPLqZ9CFCekPPdlciZt3HreaFWu5ALt81ZcxrrZRw1wLNFRktrJ1nuFSQcuTjGnuUl
8W7rwCtBr5g6ZVmNUO7jlUvYQnbvxI/v8YK7rG6SE0aKEMbtKQ+/NtfdzHGKccuwReqdDNTYoASP
7P6S0CnfgNzw/jkXNVRQg52hNHtMzRheM/GjqcZmJcQ2fHby1I7Hr4MZkUb2WkQ41IlePlXWsOOY
tNqa/3QcD+zP4vQW87+Wd0IDY4/HhS2yNt0uKOE2aoIMbgpC+I8xKGXqIiMaKaSslEhcdl+jfQLm
pdqLNH/5Oq/9sWYdbMW7WKvRROKJNMSQ7xptNeKfSChYjG1iIUxEO1Lt9+VWCT+OTgDx5gLVv9jM
FV4CVWurfO/X4p+x1a4NoUow3N1vADcSawrHaM+LLQA1HuapgihhKTHYWqOnx29TW1rG8o2TAwWH
puspfDPwYAqdKHYfL8xcR/u+MkZMMNymhDl9VepxaanWKRF0iARo/6VOK1KdvKi1Bb9ds6j1zRvc
0n6HgB7eebTqhG9ixU7qusHJ9fICdgLa5Jedt64QnrNDHKnGUGAkTJ7TO5sVRNJbdEnLYBYhyUDw
H7vMvug1WYEW+5/wtmLD4WDSdhGtGKJxltlm59ReVjfhr8XRNT1ExBNG9cZgHH9nPCnspkcQ5I/y
9LA5r0kkn/bexI9YVyp1++epfmGuSiBiMw//fRc4FRl39CeV+x9iibu+KBum54qqAMlBkcdrmLx6
XfpX2b1O3OVsmQPqBS/hdp1M4fVWZAJXp0Zd5cYTxjs0BXL3lGcrYV007jUvSWymYUEHMnpOrpmW
72whwdiq0nO89Rx7N2l4RqM/wGUers7ZOQgnmgYYo5yvcYcZlZc+Pmsa3JqMwbQWfGdqlgrrAvhk
xkS78k4jY7sBuUk/JcVWWlqozxR8Yz/+XGb8hIwO/hF3hg1WFUln8Nj52l9sGN+6lPWzO/2kosPp
YZceLjL/rneYg88Ef+IQVVNPrgVj5LVydpUPLK9bl9b5Csj36bohdBQYiEQ5AhHYKguwMs3Dc20g
qLzVjD77BNShnHo28KjVs7RkeSl4JqmJb2LosE/wvJoNEXBlw+b3eopVV5fGdf4cLp3THTyRcA9F
EOrbFtCdCQcNVitHl/0J0giZXkQGYPwAr1JSS+cZaqFAlZPpIScqEDsVuxY8A1XidccelK3Q7Wb/
mDXjcBCn+7S982eECbPJR3s/jc9niDFOGYmSWMy98AXOAqwEyMpxaiD2xUSTc5jG9Vk4U+g4AOuZ
W+8hE09kGOHEsmnscbbQ87txcHvAqFwjFPXGTJrVDgaxLSuvqg2M640kfY/UkEW32isDE6Bqdjte
O5oyOi1K/ysXRvyHxYkr8FRN7ZyLCgD8BtahoCRm/6Ik2ZAygwwMHOk5xKvzasH2mfO/UxN7VUVJ
uqNAI1ZLV4rn7C4qu8NU7U14/HjjgUtuKKYiC2YIhJTGs79HFm6mQwCo9srAcc6NvfdWgrQsulxJ
6FPrn/TSfbaU/9Ot2nlXlyUWBo2hlP4Jt5CM+QZVvVOgk12SvLlrMK8dyJziAoQ0gO8bnS2zox7z
gaj8+35or7jcLfi99A8DH5kaQvbZCJ+ncvD9QaSLg2tZa6WWb3kG6WQFgy4D0R0Zzb2wa5KSubVa
b3lA3mR526LZW0wdPt3tiXRFt1jkOr6HBeqZmtiUFdFRgU+AlMHByT481mV1rc28Q5uyuT5me3XU
fWalVHB5FnxjKjZNv6c45ulp7mFA/gbXmxt+9Yg2s8jYkATk7gNMq+1utOJzimFJxby+h+WdCB0W
ohHig8ZwW2p2rjR9y4v9ldR8OKmWdSWOMf9BRn2evfsTBTqBNNNqGVr+KQdo0Qsv9fKwk/LO/5Kd
uVlUgPwFuaAP28tsAZ+sS8kbHuSa+xEejeBvg9rrSHqtpj64720xjK3yYQEuauzCupkqI7D6FKq2
8pHb9Tl3aSngouzKA8wGeJI6GcU6Kv7Mg39S+vgS1hYE9oKgmosqEroAbDXj/mSsgfALpDA6KgiQ
iCKM07fM6KxeVY+Rpip5EqkNqrwlbVK+JMuV7R9bnfmERa/kzzgQINGWKXNVL7Nj3WmKHjH1124x
QdlSaU3A1wiOn6zS0SdGy6rJWiCfWxMrPDgvDZURn5951VqYII0dzotRIfnfFvZdgHP9SgQ6Emva
z2s2jbISY61LV4rhaDgvo21PN0Irjz6mifwrr6wnSFBYfx7K+kpEOb3a/InYj6C7xrhpv2zEQ2tt
J1RRwGF1PTMh2fInc+Z3HgV30GC3uIZ8k8xaQtkQoe4KPxk+gNUUwDw+Qk2xkwWmXjx/sINCwxQw
KyFt+MGp1qhocg5JCroADo1+d3geeYATd/RN8By+5cbQYiPZeh2dVHePmcydLhl9RZbLZQa5T+gd
u8teb+3rl0LDDuBdhpTXf+1eelO5X0hDtNNbMZh0K4Rs6jhTCSoMPLax+GR/erxRgk0774FLo+EJ
EiHwr0+KNkwbPYwHI/hYPM5Khq/4J6h4hGxAA9Q+N8UwTPn4XFeaWz6MXKQU7iyF0O5SZLk8UDv0
QQSCiEzVq253zb2YymzZCOpIROzHrzerq9xZWfcaEGT/4kqc70iEViZ2lScJaVjC2zsmMZ2iClX0
xC8WIAwI3pOgMBUfdtMW3S9XLWGKqMt2eGwYzFmBi9bQdaYl6l+LVf95LwaCPvgczapmIF3Xh+3V
mXusye00HpMLzq8d8uUJZuN7cfpogT+EtGs7FOq1pmDIGEEhBQJBczWdbyTDSygJTwj8Gt4Z/QcN
LxctDRNxtKLQSS2BpnyCYrlLAfOru81WPD6F0K7OZVSCL9wmblBIYtkY8rG87lVFviiV2j1CQex/
m2hqkJzSHKogj8HTmCAzSvwoYgYddyoiRp0qNE4EchYAx41fL22j4fY63cfvBMTLUVxqolIbC939
TlOLWyVMzBmRM72wqGJRWOqwZq9ZgjuCMYHFzKN0P0cyAXo7WsOu1CH6BCDc+5UMBKWOrdlBSC08
LiPmfXdgtCs4IYQ2WXnGRSdRwusGqNHW1uRUSXZanEQTQRdsWYnOfKzuzrYM4OjmE/ogm2YClSyy
oqsbuBxFQ7LqqmYVE+smHsOJEUbCnrjaD8vIui0IFPPI1NBPCb2spg+rdV7Cjg///Szaq+5u95ks
OdZpGDB4+kDytSLjdycLPNT1MkcnhJ3VcoVr3ykZMdner5T6ojKG8YWEeVYgB3vTiEr6UB4Zl+UG
WuW0V1HsT5fmT5aHRUCUdq71ju0Rx6IecTFLw57k91HLwBLdYv549/L0tOO1zLbKrJA/nkzjV0Uq
sHAAEPjxdDi1kB0sJ15T4oeEtDWvvOkxKaedj9UENnu+pNEETtyuO75ctNyj0Vi3Qt7lKrzyG+Yw
aggNnakZLe3LknjLUzslCiyGzUh6F25iI8rFj9CJiP3JIEolybl8AaHXEqdZxx+owm4/fnMY8RzI
kiDDrh2oFwavwMXHQlTMF2fr82jTHqgvCxta1Yauavkl6i/IQP7JQVSPfDRNEojdbc0GOTOTjoO0
PNFp2+TkjNfI8qxxmE5Kcw7AdjEMaVRldZx3rxe02H3IqUR4guic45VDayIPeOsvOmDZg4lwJTws
m87ksBCYHpWx4bPavCn4/pcDgojP8Y84mfsjTF3NF3v05k6V0eoenz9dHw0ITFv9iXGzmLEmGMK9
NOTo1jTFerMwj7MgnmtBIVYUCwtaPx3YYXpSbAC3vlWM6scE8IZJniL8E+bpCKLXFnHt8p98hyZh
kfeoIgArEXBw3VVTj3SjAhE7acE/JLLyabFNl5fXOaOKfOkB0LRjPQ16FKBLxztx4MsznFvJNZv1
lA7Y0jFPyiKg530uQeRqNyGz5rAT1Q7XkJTHeHWuCOzfwHV3oYV94rn/+kBVsSvQr5l+eI33YRrF
196nsRD5eGs76zqIzZxnBotKczc+uAysxRWDuabte+gnwAMGpKBHAO5BygR5vK54C2RDxN0lh7d2
8bQln6uIjE2X64B055q3ZN7JG0GIv4yptygKsIyrwMNCGLMPfl3L1N4iTC1c1sZOadyE+Z2G05IV
LpgixGOBUMrsuw5wwgUc+pdEF6hyIXhYlNCcraThTra3/fGMZjXvJZsZfkUKlH8z37Qv+npmmkWn
UOFErF+Z49ilB76UDu77qyd06uNjcNeSqbgZSpFBdK1IUHxmi8v2a3U3Ll0DtcEMUa7dg18/z6Yh
xSO93TV3vrljDKq4qp9/QCpTGMLmE/zcQ5Fdz9RqeHchtMLfKHeO2oaxFS1/hG4DdSckrzf1u0Ik
T3bsfk6v5uGjVar+r7FFJHuvGv525GZMOMFwYz8DQS/suCuGamM6MBWdwxb1glIZvqvVA2vlk3c1
ML2uHw182Ek6MVr+T80MNeoMg8gePta6cNu3kt8dqKMuUhyJrXttkHGzBZsjlP6Kjfu3LV5LPqLA
2n3FI+wZjC6iI6co6zNyVka3DDCjrwOst5e2hVPqCJE7IpIkMAa4JrmcG89vcDr8OfQMNc+Q60iR
rVt+Em6x62o9q7dtzqar9cae4cjbougw7XZYhT8Z/DXCfkWhnhWANtgT+vgxNgtsyqra9V9nRY49
EQsqFC102/g5uXYh9HawRmOA/A2lu7cxHuJpq+OBabG/4ZiwyzXdB1kxa3bzUmPzrwLUjGWDOgJF
tW5uAX3RVhElCdMmbWvIdQ0pZf1rIStkQ52NZhsjzk978dNzJ2NxX2lQGQgNkqWMLTdFvoA7/jb+
lz14V/1lQBDr3IUae76NVzxciMyCwdtrQBS4ZcvfkF2MDBvmsyhc9xXfgLSjzsejAdcMNNyMRt1g
bkHn/SxLsp2JdSj7rMcAk3/PJS8ceDPSz6A2qkDlVNFlIly3vEMUwXkMUfL65NP3hjjXRLXw9mjO
MTP6aZDsNfuFP59U+ogwfTOrACXy1HaoBIUt2BohUwwig7E10x+XRfuDgBfCezOevM+pAkWxje3T
Tz6/PS5zDXzsamBACgt6SFct4dj+MUecvuzQw8siK+0t8kunVd4r3VXY6CTizK7ys1XOgrKzLmE2
pyggURwQLsOi9Xc8CUI9JsXnY71FIfH1VznoOJcnqp+tx/40FK8wQZQkD1iQz/hIKxr1PWZp55t4
KKdYaVB408OkKl0Jpxl+4aRNCs+xv4P+sKyeRhi8qjBI5YVziJNpSoPxsFlDe1eZekzLKcNbIMK3
hdZlL3RVAq3jIWkmh8DZfOM2Dbaw+h8Gi8ictWkUYW/1TFVXHnC9WpCxCcKfpR+9WS50+j4hUsZO
PaNiwmE0LXYH0B4mq5N23M+JsFEyIG/ISkRVRgtSfn/y79fOPYWIEeXs1UoILS/y+0p7MRmjfG86
vo5d1BXgURGY4rScUo3FJLv5YfVnAtdO+wpCU5U9LIcBo2kFaA2PGTU/W7d7TDIyfgJquc5CMTeH
aBDP0vTQcFH76wSEjOUJkCTbs/Es1zczZgKmD/o91qMQs3WuZZXlNUx7xEERWzDs891UloSk3RAU
ifDqmR2wEbHvT6FWRLerJb2gQ8XDzgHyfS/TW2vep4I74mWu9OBOl68Cozx1uOgg6M8wUhfpvab2
wqWg53goUVmZQtxQKYQ0aJjf7tbHVYF6XKfOeG68W5ghaMzS1g6Q9cx3XarazRRpAaVk8Q+LYNJJ
y1qfxlkuFJeovU4Sj8FMH3eF4Z+VQaqQRRIq4/kSRW5uZOEZOjdZt3eE4sP86HqZCVkYNL3OUeub
nvJQHTYttCSFL3WbGBoltarA+X3S/6bH783XHUC78+C6I/Qx77P3uPnecRdGRFh6VIstu7/YsPUz
3o9x/4XoUGokUBlZmUFb7HTINZrKorcvVXHSmNmEqPP7i5QDDWdi/jUHRtoq1gZm3xfZEtAQtWJr
kdVasMWsjoy+8/Yc6zlY8jReD2JYEOwph0mf0TD7El/htVetaGtZ6Wo1mZ+BFdoiKuEm0+0hNYp5
tjqhkhzT8w8PvsKDaDWMtvqi3w/OhYg0wi4WVj9bETLvXk3/TNrLQcsE7NaNpeJWTxGWvLMINiOb
t0v6TtKqaAFT1emgfrQIuj8PRcTNIUFcIsHozXKsPsP3F/JxFIZm5QEBCoA1abmMXRP8jcvEYiEY
76wdVoY28cKPapXWHPbl7GtkGFizLpBtoYhq/Z+GH1yCjlRgmsbVssXypRB9JBGJRAL+02peJ8+H
7F1+pxVWPljcPeBt7dFBSPX00abjOXNg/WFSp3rSrKgHYamohZV2L0Gn6Eg7Ura7pJ5rrdtkkiUW
KGqd+jEVKuqb0AHjCEN0fYZERBvdmLSBO/k4HYYVGYi3j9yBTXyvMR2XlFntHHT302vIcokRz9rg
gN/mGa9YRLxOi1Ek9lI0WBGH/xd9XXWdwFjJ+iq2FuKW5xn5rA+VJik+FWiHU3H5uRN/PyO0FjON
m6ZMuLSWzQDiccJvj5jPc2g3z3W8n78xXtcbblk9Vb4RmYLS9L/IHcuFRqeM0fXTBp1rsOIyC5nJ
I5AXvqBWvWIq2C2MejU0VbZsOfxgW8RIxBIPutW2szOzzQPueby2lMqlcwSN4iG5n0xxSX9T+zjm
33D/DcEo+DPUuVL+/lKeGPLKg+0x7/MVC2nKX4DYhomVObiRZ9LAf/5Vwx8+ODBjGD2mYJcKdFJF
BiHEBHp/ZKaGZev7QFOqsqcgJkOCmsnXX9vFLbVLLRUDY72EvoKRB9HRzaDJNqsnSFIgQVB8Qljz
hlSPDYoUPsng6MXxGi32UsHzSBNvV4GbMzah5IFIdvQPLRUyr08TZ2mcXGgXIu0pyLjIkTNwSWoK
4pdKj5xUx9H+lUZqZL434B1rm2VcC9AfeQ1S8JSOGU2v9K7wEMw1djIGFsIRovgXZ6Fu/jrcq6OF
vDKdCZdR4RVS6zSej2p8u1GJrV3VRKmL8qczeCjND+wNG9zNzpqvROxXQiHfoVVxhnqzFwYBfhDg
wPbrM6zY4rzd5eLI1HKSOpHFLAVSvsKylEOejvWGMKYnt6BV6XiMNwGa2OkxNkKFF1hPaVqj/5xM
9ftm0GJq5JOHb1lOIK7byFR4lZlwHRLcENlrV0H+9vq5wspWeSdaMzxULUxZM4+RbN99zbHXsUb6
UepomVTDJt7j16xE94MR9sEP5jAm8uGBbmqnKKKc5YYC4YXAkZA5aPBcayXn1sU/Tg4YwmpRVTMu
NOgNWR7lTAL2qbUQPMQKqGyCXPkGLK7o8Q402ZRL7r6VkWFfnXTPK1hsyTy8LzBi2eCdY2RMeDeo
KeVneymGKdfg6jFPndZY3lquDMhBAB08StvHPxQ4Poi/HRJ22j0XV55BaDArV/lD+j0wc052Xddp
qrFgQpZaGKebIB5t9iUthYh6DuIKdeE+8wu3EihcMTV9B0Ce5LtgBcEeiSyIACRN+QK9z0oqUbg8
NKSg+Kd/xcsLIEYzsUaadodWkTOUtiBgrPcB3ZiBUoemIsS5igDuWI6TMKcn9BSi7xVz3IOGFJA8
V/mR6PX/Ii30GLCprTZjpD/V2VGkWpcZva1WmWBVfVolCKf5KPHttieAL1VqG4VwnAo89P/8fOrc
XJvPp3NagDB3Xc/rta3J0dAfT4z8iA0F0ByDClsOttAxa9mWCWrOFAw6z2vBLrBVKUY5mUDXsdLZ
MQs487nOuVM20u44eqFtEl6j63LKqGBgWATE/Ne7MkZd/mdibTiX5x9O4ZzAH1jk/kr5lVIvyL8C
LwmwCq2XUIQsPRqbN8TGDuenlifQFd0KSXpsFWumMG13fJmY3TTdmbXxHvJ4EVmIid1044mK0oDK
cc2MB6bih3NRPAbjP/46y4ZHqoy0behzWZTvXTKKJuqBaWyV9YOeJErmQJxXB8FOPqWO6voik+Ti
MVlT4gRhHoozL5sf3kMAzyT4oxDXQuDmXXmL/l3IsZ83LSI154RR7danPnqM9jsL+Uawa+1uPuoc
VmFngOV6hfLv2zzLsyGuSlba2/AgyGD6I0ry5H4MKYTw3t1DzdROn21Pf+8YDBpCAlJzcEd2WvBG
spAQy5ilznQ5PXgwThJDXVALfBOZJRR8yaCaEXkHs8qOmt22Ox6wy/dqLpdAqaJhJpbek+dzRIaa
ApBqGhD3R665ecoftc9fz27Bqw6CuEWQTBWLYWTrF66FsNI1RmMdtDR2aJOafjKo/spIRHDea0zo
geXhC9A266JM7HCuctaXDeCt2aGgrKvypbn4qy4RB33IKyzWjImaqEaEcTn2mSoGI04lkX6VbGy1
+aomW49vb0L56W99SEX+XvPCkc3dKRcKgRhdIKJTaU3YYdNnxYUKLitRgBBODafhrgW0Mt+mLSMa
vcyFIyAGpPJY5+92mIykTcTuF+llrFAPFpRPYl8bBrekwrXMyNEtlFIqA7VzBSPisK8Wi4763kO0
jebz/Zo+W/TbbhW+A42+VvPpzGYoRq7WBn5jdynebo48dqLaslUKgv26p2qeD5WJyHc7wQ+xF7t2
N3igoApzGeTuEIdFYkuViE/Wc1seBsze7WeySbEd1C2XEn7YTae4vfWq0VdQzZVvS5aZb1SjkQuK
HlJTuSb+ZDPCmMnYC4DHCt6swuy9Jm0XQV2FysuGZ6uT1AcVLiE6ZomKIJzx9HYp6yokLGI1RaU+
Ltlx6edweHatMb3whJRtRhI2UajTGeUdhftyOebulnvHNDoNvm2eEiCatrFVUUDU/o8bNn3EE+wW
+H59TnPs0LhvkBlaY0Jvv1WBWsllV7q/fnvuNsNPpkRyWrig0LBEzgBrGpKaGJB6ljglG6YWgDZL
Dtm9xOL37tD3iteVnLh1BsMpGIiYQwzzAP7gIw4oY1PIwtob9RPn+3b24sdRthwy3Q0ayyog1t2y
bx9NNXXWc6ND30uDs5UGFUYaUVciR043sCN1pFdxOIcfdj/pDGbZqEu9w/aGz1abPF7fn97xlzrS
kiN4Vs7U5Z9SCcBEuNV6P0apRneodX5V2icwZZ+6quGzUUc5cYkkjGpzI4mVCk/uFn82EmMrFPk3
udt2sOtHcvsoIAQbi+cRrHADxQgQVeOA/dMXYxQqq7FC+ulARTHFQAPQN1iPxLw4LhVgY/n2qmB4
weYhMrnpPiM3X9lXMBgYebcaHBfdkYtDJJIMcjQe9FzdDcW71RjnP9bbmdfGDFwWnjLE+eITHux2
IbrIOeBuWkY7uN0gQr0oOb+/2zPc1X1lG0HSXVwZfoLih7ZvdhCqlu5xoDuxGt8ZgCrN1wDAWmpi
1i/ZhwmwVbDBpC8ggXY9L7k/P/eRObr24kEA2lmWD9zSH+yXMQOiDHhEXvgqXgmzHTKaR09mIu5Q
50jiQST3/juac3uJkvHbWMP34UnjJlokHjOB6hjG7aa8o6uEs9aKeaWvkdFO6HTJqfHlhVKM33yy
rkzPU6x80hpwNFH91iQNMFC/0ewipE60HmGWwVcQSvWiU5SyOhs2ATS1KS1b5DAiNgTzFV+Y+RE7
QszCd91TVGHCNKwdM9eKyCLJAzaQe2SWAmyuEy1VWsswoCiOJzMfuYYkfO43kG1+87NRVSnxKQyz
SabE1EAPHObSi9rUGSGi/b4i/rcnv/45927KJ7SzV78Xh/I7yVN1SuZI7zaGCa0mMZX4Ba5cfBwn
DHjRGT0uUDwsfmoF6akY415U0Kn+vcAvl2Rvf14e/MKeQlJb17W5dF+KmEn5juuyYS4ncwvvwtxS
PL43uVwCW1gdXgbA3CB2tuLFvKXt1dyQzt+rwkWD9yw5ZUkwS30GMEjBWIEsoEUmMyd21PkXtEIN
zhzolb1zmZao7bnmdstn4hG8uJFIO9LIb4Bsv620cVoL3k/geIE3tloiFd6fovNk+84dOQYHsIUn
RBx+Mq4nDyskzgyQBl8CMHJkOHPJYlKgihdXac7sfahgZVHPkIIZXeTOHgQ6A9HQo7ioP0G34sZ1
DAE5F5/GP2xEmgsj5QT9xra7vCE441lPCL0CgZuENx63v1JByUbQv3cPmv94fx6wplTWPgTQ/MHb
lTHfuHQtkf2U3NzOlFgcSc7U5TgvvrzKWtPZkaKWTeExyuQgTH+MZwozHldXJKsR4OGGWLTCBpFe
RAXu2Wt3F7sKXfFq9I81xck71HzL2q909/+jZzvOFUKvzm7TcTvMcgASOT4k+3uLXa15hJmKj2p3
KZrivsVvHWreT7MOTCZq48UdJutbGtq4/w0Uffjxp+lGxCfSL9pxD8LIeoaDuJIP+Drg/bNAos2f
ri7WzY5NfvFywn2RNdwZGXVhFx51Izvtxa2TMOjJTCW0uvIr4HDiG43wIlzNw+BReNqvOty9bJRk
dXrxuY+wVKCiGgl7f/4RGiF5+fvM+1AuQPAvHq+7WWEw6hEabeQwUMY1+4H8Y7S2bfhggJ5NJrzW
2TzbJAvRv4A0T1y44k0f12WgIT1bnLyrhJCWxmru5qyOHqvIPFrLS+OT/fGQuTqnMxb9zw4k4PCb
/p8pod4CTqRd+0zTsMdxuU0xjqEdaKXrBYjqU7iDLY009uZWNZlkvhC/tq8q1o3pK3yjY3A5keUK
S3mS1guZsG6jvUkqncIcj74Xs+txOks7N+SFsq/APXef4/EE9Y+4u0C9zQr4zRjjNpG/QFyoWA/E
Hba5CvpI8CNQn9xjAj04Tc/ynuYmmYziDKzNSul+GQifRnvoQonWAI5Yp4FaE9eB5khGH/DrXg8I
oz+PqrivKptdJPBQgcDkQducQ3zPPZsLh0uPm3VXxs9h9OHIzZ6lkArj5nionkgNho4d1gCQNxnG
u5f96zUIUtlkSUDzWiGsCs4gOSpvZIqegXRyzAXfQk5mEdYuLWjcORl+ezc1g5o/ERgcRgNtmvuP
/A6jXNLxn+W9ONodw1r3CHeYxYMVLRnjsimS2g0TRIAqM1GXqR3vzMXUIJqsig1k+M+BvtSDlSyK
KP7z9o7TdePKeiCOTca/6Gp0Z3zPRfnxwBILolkJXeDkd7ecH85YwGA232Pz1lTwjJtdgPSpeAp6
LxzeteNZjWLXJQxbM7JKipQml8m2wWfQeDVf+mqKeiOJV+Z9mhgKniaKvaQTJjta34pEhhp9flff
YhMS/+ksvr6FtbCp8G7j4q+niMvRK51vhNmk9mwyK50UF60Y2+VcJaldYQT9PGdmMFR36CHEZGkF
cZzf1pntGQG2oK3UXtRp1zGy3cJNbWt26cEuTNPvuiARXHAY8TK2jpf4D8SDIwgwo6WmSMk8jkv2
EuxtKZxqMrKeCSKxyOk6yjHwkSEFPXka2KKjuX4kreAgR9bjKpORFgNQ+tRFgEC7rHa0BlAH3HXk
bp0IQ6PeWKBRwD3KnoyaqH/NJnHTxrWtPKZUzW0gHNKSdcRCDBGE547BPD7rq36HbVZ6IGZkaBaD
yGpMzY2swhPF3OEZa+DmNUV0c0Wv69VbAMI1aw92MOO3JMVUYhKtink8lwVVe3Vx6cg9l17bbpMH
EZGICgZw9NuCuunfjLjVuCkY87ZcHZSqzmsl/epsqYmvSJmMTsM9NosqI0CEV42bXlGy5Z2ef55S
GPbQyAZNnr+QWasbMyg3gzcMnF0zG4Pz/WG1gN3vQjUlPkp3u3BqGGohyd53BpBoNMZADH1xA0kL
XkD/p7nw2xBzlEPfmi5led58aYeaeXovz7Gkfoe3d74s3lmj0VD+GSGp5CMXe5s31/eWCzqKab5O
+LiHTMSBF4kRMsGkIu1K7TZR5O94Mpo7ABBz4OV+ox06P9ru9XM1lqtfaSQt0IB+PD/OCfeYsLeu
D1MBVJMfG4wFEWOLtT30s6QtCJxObgThd1YkM4vfrohdYdT7dea6UeE0/NO0+UrOv0xCOLC5TIPk
yWrDR/3xhE9lur63AHxJj4BU3CvgEGngesrcdbqVRcKOrU7Azr7Aq6Unrnx/hCt6AfoXNmfe3VsG
gHkpyULBlzgNxqFM5OyKbYOEbRE8n7uUUDx+YT7Kol05OfWIJbjbLqqRXpN9Su9djj/9WhJpOLu7
URtQ/QUdFm6knxb4FudhvW6r9Xx4lKWG+64vkeVID7yNWh68VpJxVzy6zkfBvubHz5m0OR7P9v4W
kGuIhdQC7cXRWDwPIdpHO9xMkqNWtjRmNSOXqHN5uC2VBGnx9C+4hhnrMPfhIJa7Suq/zlZmNgWp
5heZXLWCWQZPa6c6ZDV5/5450t4SQfCeCoxa+9SGClUwoyIKqQfk8pK6Ht3GBBTTYcOdzLrGEauE
Vmext7CI2YzMi8SJJQVOlOWk/aYeWe1j3PRpr10MrUoEsqUm/Y2BNn4IXVhTLFvxqv6eChBmQniG
2cNJEXmJcRmvO8ynXDT/aBQF3nsaYW54u98u126l8C/BNImlO+aSW7bJyZLMRixHkjhuFLTeKK/p
iViTBLXQjiPg7IJCIZp7YZOOvVk6blzz6KzPcdx7ypXMUeEUkgzJybcpVA+ssHidN7swgC686aGh
aUrLxnLlZXoNJ0fjFRjfS0/w/jGp5CTipUMdW19sVyaLFewnVRGPFRh5qGp25a2K+2NzPSNaiW3e
szZNN+cjpeu54VtRmYfG9PB9pLiH2TQZvWu2NU7uMn3+UvE2q+J1vh0bOLZ+LmZIbMY7MTZ2+Mme
2tCCvnYe1YV9SJaBi4qOGg/W1l0Bqw48GqgPDq8yB7QDC76CyEEXimldROZUCTlYmjgbBPyNBhZo
YcU3e0itE9rO7BZ4yCL/hrQlI5x13v9nseLsXtCq6J8XM/yLfjxIbxEXGCr5jerAuneOUvOcQfOk
Hj2JoSGl0UBfT8m1YHWwUUVc4zbkF2rRPMNGFuvXxcCBd6GCO4sznUOp0K9trpNMqjRKq0ooOTxs
AZUYOOsGQmPypWSCwPzuJMxQvq1EmS3Jq9rH7NbwmhqIZSvK1OL/wnbAm44JacJ8Ed+oBV0OMzoz
TNlvWgoE2o8b35I2SaDeayNUaQRV2kQTR3zYnPtnCD7v9WKpZ7+gXYWITTkg3Ldcbw6WUBCM6l2g
90vVB5jnD3gf5fw9z/UFkbYFBcT1NMMboj5mjm+tj3R6ndOx03IUizY5h67HDaZtKqvhtgBt3Mjv
YFbCcpexa9treyPJtTeM2o/Get4jd75vCRT7hRMTM9O90vsxesFu6HJtO1y/h9rxWs6C1GTtD75C
RMnPF5JYgrBjXhjD+QQcOKzYTVnBbNfg29HVzKu0NKNYczaxxVtMLkDScJgDExHoWhkZc0phpRIJ
3wW0p0SLGGuImjIgv3EOJwCNoKM7t1OIFAlzXpAp1lv/mDu03gBc9b4yHSCFRWmEgRCdeLA5K9GT
/mB77oNhPATF8mTSXs7ka+jGTITiXsGReHrHDVQtWPgOrOeKGQjfU15xNQRfIrKl1loUzMfxpsS9
BFxj8AKFCkjQgbBCCXehYOHk8ylIfpKwFtZGEZNvJWwNRai6tOOc8Alsul1pcyw3sai2SajzGxi1
UnOtjV3aSpSIsIcQkHHUxHbnaxe1dBthqIB9MpPVrM4DtloLXMZIb63E3WrOfFq4OkmgS6a+VDPi
rElnx4aYTwDyQxvcD7tjB5rVnH/ObSKdhRoazXtQZ8jgNPXL7uKiunxI1vXTb/C9eRLv8xuyQQN0
fSyrTobkIWqG73ZqyMC7TE7XwBsDSCuLUiX1GGr2EN+OD9kCYgam21gQxBM8Nljt/+buh4N5egPd
irtHYBC3uLf7cUTDeNOSgqOFucX9K6Y5ujCGLrtbiZme0O3GBrHPuIMe486N94PFTaqCKk2PmzTY
2Im5wwJYWvRjoq+FlSmaRKrwYhA2r/Z6JRwk8AZKVfvYRzV8sFf7NNliUtSZokRgHicHOsFYMFMj
iD6kx/8zQKpWGxTM0NZzYMF0dei7V86Cq9k9YK0Igf7JaKifA5e5oHnKpwKyg1AMy64IlpdalGuI
zl6hlED0a0cgunBzuA9WWddM3oMpAAyjwDAmijw411nzUIjoMSbixWlMtu9rYzwYjmK4VRkssINx
fgntscAZ1j3iT51/lR6ukI7Q3PfcsvSC7+obX/fM+Q+4QayOXrIzxzcplUbnYOYfURLN7FnHRP1u
DPtCL1RnO7EIFH5lqtwnrmcona1kBTeKIxes/y788rYPpTjhtXYhZk5NwD2d8hEWorqS7VXFIeq4
hWscLZwRpRl78qQN9WIN0fZauOXAupPNkwkLheI441j6rAl2G71C5mz2GZ2H9nPYvpJeaIMRx8Xs
m9IHj39zya+mNcomIGPqfJpz5yKa7ZJLXXiaayLS8AIcj0QYlzDF+fUMSbPfsWvreaxCBOu/e294
et0kpm4tl28VKfAfmCNQYtfrSHENEghrzfLo6M4VyXB31fVG9MUuc+QPtL1AI22ZYW6bNrK1ChTs
KpsFsVywbkZmAAGS6gBEcFZbPdrtRu7sSh1eqAuytSTVA4xeWxcMumXedvbR46j/u6xqdqdScmE5
OdNtksBLhVddaucIfI8kVZO3KXWyRtDiSVi28NXmv+zCgD0UzXjgSQ4IIxYGu01uyuoVpRAnoH35
6cr2K/QDCLk/yx/8Q8KM+wYF2XFK7pop7Rlkvx8o2Jyfe7W4OHTvTBi2nkByVK5yHLLu7XFHFFq4
NRHd5OJTfSnceOiYnjUlAu7eEZC64/LkUw6bCeX3X+phM0SKbR0iMnbZO5o/oe22/LF943F22jAs
uVQ906orJI6cAjn4zqwmoOEy5Su3QM97hyvURLbQrlA++sFZiwci5XfkY+JKWLfmxCFH9tazVU4E
kunZv31twHmVhgFQ45NSQ63lIHgSPcjkxWaPjcwPb9/VlV16seE/ju6u3uw4IEFvdC3QNqf2SKqI
NhNk7bo8Ql8TUKiCCb5LT1Sbm86UiFvu+h/R8Hq9SS5ZzQVPlwD/+v/8Z4AfE8ForfPDXlCzqOd2
ap6S1NQJrNgXwXvx8BfDzN9pIoe9KKiEbq75CW1DSg20D1NZCJbK+4aEWKhN6XtuLwPor5KUcHV0
Am0YmPjB/56QRP1TNIdlqMtK+X7b8bEJFYd80AhSzoBlhG5qPPibQJgrW/hGsjO4uHGdkRgF2xXk
BenPLPhuhk/28tGrOMRt8ybw4RfqpLLVcwl9908RHOOsu/+32ukc4zKgoiz6GbsVGzZUbSDx1iWR
1/tA0BnnZf75ennv4oJcCb47iId1r6Mf4ghr1vooVF3V+DSLEDpliNWYb8omrj6R3bJ4TTT2Sxsr
NvUUzrCDHILparwAkEXcs6+UuURlQ5Ur5hrkM6dwG1+cchpZQx3yvYo31w82exGhBNq71Imu01HI
N29g9E/qzs4NUICTlNgHnTosbT4FkaCfoshn0CzKBrv82lz95nv3ohASQpYEvQKCTUx/Iz0bsN5I
MKvaPPoDsBtCYwH8jX2e13yH83suwrgDK7UIGhIKLpWWHttjUKB7zFA+4ICpBM7Iw3mqJhGVUDqe
kxNvd9otnLxrrI/+A9qfbcZxe3cYcQIC2n86NloOkQ+LhMXK90KDRmt6j+YT1YTA1voxvZKBb2+J
SCsL7DUExbV7+gKfWqjiZWTNGije9JM0bU8SeaRC5mMkShAQkED4aajnbwPw4Aj/eQ5Kse+u87Y5
5ehsqc+8ypE5jUHolkDQFUioPliOILRzSOJGbLQif1BDGydS9woa4XNW6UGMp4oUwmZE/0nK++Qb
t+ua4wfmDSyUoca4s4OSuIp7fl94700jtbbZn/jx3dAachChvmRaiB7Tgejxz07EuTuB2UDcBpKB
XdsSlrVMZzJaWbX/MFf18Ur2Z/i6hr/e6mNy+rke1C/+vwdqRpWRtv8XOa6EEdWmkldBf4U+NRe4
BRcmluho2vDaeYw3AeLfLCaVrbRqdKBEAJtrAJvCTCouR/SIvleyPNGA/Oh1Xv3BBJJrNr4e8KT1
X4xpqTiOBq6jLBfhJzvnY6GXCv2iMP9jQ2o+CT/HxCDOJcv4jagtTWwdp1PW4ceftkkOAopi2VSV
plKg6DqfrZnNX5Jn9fslFJwhZUXa60UJFv41aVxBI9BkOmO/wTAjtGuLXseqaHaFG7vcoHnYKbju
deCxb+qbGxgzIUaEc3Za3wzjq+b0oG80rVrmDiu5jYOUsooc/WsBqXxTL+beywYbrwWHbpaceZot
jdKuInTKMpZBdDdGP/1dcQuGeLUQrpCSujX3PAjPxiy3WZ7wABQk5DUtf9B07IRm4yUMeBf7t9bp
/PQGD4mK62WojtCaplEo13JzkO1I9NPdRnWvOzJC54mgukm5WI3TPyGZ8fO2S36KMfCWRq4CbzEZ
fZ9qaPf5bqOocI2CCrm+hfK+9GuWM+CEoqnCcWmSKgiY3Eq0kiAhgEbAfuwubB+GHlWjC+6m46fK
toE2V3ixRWx+TqmiLq3CI4i2FXAiYd3V04OAbEd4Z8UoR0fwTERnssRTGag9tk7d2tTlgkp6HzGt
iWBzR/bgy+muXqbNQEHZ177oTH7gKEWpLwZgYg06yf6APbAq1K5OBkZ/5Nhk/mvUwhlNxmkRqEQY
1IxOaX6Pv2LbxAPQKj6pH8DtGIay5LXsDIR6SgymPVL0/e67HKQGOuIMZAcF2OazuU8yNgklO+pw
hc73o0xx0m9Xbq1QyegRiNhb7fLsoHFGkQXGbLItdEmBswZVCVgn0lkuQbo4cnlZ8WpShrTYpHqa
lEc02px0vv6iLVGsXP7KV+r3ff/VLdDQgeH7ODGDjUEy9KN+5cZBkJEDA8f2hvtMIrGYkA+V54Uw
redMNX43D52LR4Q4wY+OmEVg4vfzcYiD6APIURXQPKdUVjNDn5JbLQcf/UXdMD/BYVWeZ29d/dBE
K3Um2U12TppfeE7VnQlxrSqHhGdtUzOUE2aNpYD8LnX/BHK09dIBYr6Ry/kcpKxWZtFBWBqOHQu3
Wc5XXDzoKc9ZF8ACWtWe6upVJ1am/Zt9BR9K3uAf7lE0rdke1CiAqnrKTIf68hoDJ+pUuXfQld2i
PPbqgQIVDhLxOnH6U9KvXRHfGRsVQjzLu6MYalK8wAGB/3jQFmVxdjvcRFg3Ms8ba3qvIALlAN76
SbmktmhsmFUoKrW7/EeWKyAvuII52IQnRVVruFLYQrvcCNHytwIF+oV3im56F71EdHIehJG+Qe36
s0PYIvQKm3zU4UniK4T4RpKFM/QXDZkhz1qZI7orMC/9+tV1L+ultCAOi6zTlQztIv4fhkpy0det
ytVdP4nOrBMg1aotVWkFz+OouxKkYUQrREMHUeVair9CbVo5oBpHOf2GGXe2JkylIhEm48VyBTtR
L/h5F277r9fd+w3vPD8t4s1FG4/5Wx21NcWr3fFvkGNe+TL/ml8Zb7FR+/dY22WUtX2uD8zprWs6
pV5F/62GbPVcoZLy4hfWiiwQR3MBAk4yxmD0lg33DoTDg9gtE0u7JpYNERxNMYL/6zN/alf5b6X6
URMuTRdhMkY7SIJs59iNMwSaNBHPUi82N6oq4v6wSXDWKyUcEfAgh/QklklFLehB5pBI9HjmXLZ9
mfKMRjWb5GTeftGLLnPjw0clCgvgsF1TFWENtwff7+aJm5S9vNTdFTck6k37gQm4vIPF0QJXVwM/
UGJA7eBFj2+BJD3USN2KOtWgxspe14+d72GQjdbVTbj2uLWnyktD2jKmwIKeKYrN1nryKWzMAprb
zldbPKLQc2PcRmD/q8sonqfOFwn+LiE3AvPzQXhBnACu5I7PyGzyd2r/0xT/kbvr4leD/Ts8n6Gq
Dks2mQ38Zs0bLi8c5QTKFFe+qEHLNxOq30b2E7vmdnZwBd5UrfTU1XLo14SgkYV0TyMWAVxD5UC4
+rMB5NL9zYNaapCH1ixB6kja8DJ9glFtBPve05S0N2sVNE3k7Cd8IUZbfb0bYfBTCMfZBjrpbJB3
X03RdL83RXEC9EFkKq0FFowLt+KNt9vVQvgx1tNQsmqjjSurAwdWY+BK1d1ve7OrpbT2/VeOlW77
Ywl40EX4HT4VyNP23oLjPaC4zStL2ldVcIcdCzr3SazppmPaE1b2LUjVleBQRKNPV7WRVV4YdGzH
QOlZqiV9SWWU/X3+9WVy5B6e8NjAtrPhhzT1QhafYtJjvWimDykU55R55TuPW6l3aQELunugejRU
l/Nnicxnd4o2x9OdKmRLlVca8xMeeAfVZ9IgZGALPLgixYfQFI/ARh8jHWiEHxJ9XxMwbJXWPniV
qzXheP9rXVHaU2aV3P/lFZOj8NGRAH194T6wYHNnwpRDFhGmREQM3bK9/yFmcxtr/CGO7vqL4Syf
8p4VFlVLxtdEpzch/g6KHuHEVfswZu21DdhNTM1f0zNKY9zhXh7DnA6aYVtVfsZYz8i/2v18nCwv
fSA69EvHDc4bNvqf/MbLW2SgU9jgZAg+7kgzK1xeSLG2mInxKKknGPW8OQ7CuLEpjmFjJnLE1Raf
L1jTiJ9JF7BT+NNKh1Gh65hSslVD6/wALZywJEch6v6fghQcwOKn6hbLQvVH6u0i2Z95ERITwxnl
j8sVUwK8yBDvm7iubXDHZNS3CPelDndl8ZRXBewcI3dv4vkf92jBVpMuSs+t5Zo0DXkn7IRt6M//
81DDMW4Eb5HeNxTws9n6uX6wMZ/syLOEJvl/8NCdcGdLv05ecxh/+soShb8eiNsKLH67OpDBAI25
Z4PebOUexgVbSZgTdvrtG1as+RI52EXrQDk1DO6hu1i/Y9HVQ4Gpg2LHa50sdk63jWMzYmFUwoYH
ETkA96hHYpxqP48a916AFtSDXhn4QetQFv0gZQjkK2gbiw/+7un3KNE1L6rr9ltQZXdQpG+jasfL
V995K68gVTyB7mtTu/1l7RmJf/alsh5bBBppGE0iYxZ/qi3hg4TwMiV2jTNBOnQ+7DscowRUnafQ
b5nCQsFBVr22rGnekz48Xj4IJNZpNArvnnbv4sF8B/z+JyAEEUKo+PRMFS6H1ugjxbKeI5TP3+8M
SLztHlZstRjogJv3kiY6mKolDDZ2jc/y+8N+RrQDvikz60yCcNqZsncpWCyHVfDqVancqfpOVQU6
3xow9gRa70eX5PHkEi95VL5ovXtY29GwHxXZOMzjh2L7vd0F2gMZGQwMUA1QCWaHTRzCajfB/016
LwNQAwF0/3wJolfWhcDXC9iVe1cng0P+hAkjzvg2hHCjMSRH0pyOFWPI6T1yWlGhJ2CzqOP90u51
s5m3PfR/Bo/nugUzzYyuacZ0VCasqLP4JXp5D1ygweOzhiwhze9+eVjcg4HhBnergdbPbzuc9H4m
ChZYIHRrvoea7GFfVp/f6LRG4i6nYwSwQqpMZV7gC/23TYn+Ums7qZi7zYDmNg7iVX17qtiRADOz
MAOQZerIBTbosu27+Bx0R2d4rKodTqrLPkM25Wt+3IpTee9FPZLvuQN0X7b8HvR7HDnlTCafyiAt
BYQQUh2Ygg3XpY4XPnsxZfc7M1IVZT5+vfO8CZnGUAZvcKwhGzPm3kiP43fQkLlq1kjd/G4Wp2vl
/fiZR/FMpSJlf1/wCRLT7lszyBfTv/Gpb4jjay00HMte5MT729wyl8EMsLs3UXQYII1hTFjZUZqE
Tdjo2iLT7iOPSVJ1xH/MpBWnVGCVJd1QIhG12TvTtCR3LQlVi5r+W08tELMMDjQzwb62l98PzbMg
gEZU8HoF25u8N2inDak8UBVouklvVtdaxGAAK7jZUu3rw0kPi6NK81KLL5MCfNmtQm5Uo1rLiVb1
ftwk5EhO/kMTb5TYjiLF7S/1YzYJLtj897iV52pYO84UhZl5IOtoSZ56BCItf6CSOdwDJqkTowDg
Ez2kSdQhkUbQoWK6kjxAkom8GOkLn6uzveOhfD3TDx0dlYDBABdd/ZtBdECwuc+QUcYREIJ29ztV
VGcM+uGSV7fJAA+YIxBJzqnwPLp0O155NZe9mWVs9i9yjs2l0tipnWTgMJIAwRRnIqb+0jPgzYbw
YatGcyxpKkkC3tza7GEE2hBnk6INy+OqoR9ON5SB6EPUqQZ9KF4OP2ZrYr7nhrf+F8Xy9zTDbUoP
pCg3GFi2teo/pid5kBYo0Y7uFfd/IG23KKUmlHJ4j8rUFq5/iPZcbu7j16/ADEmG9yAJBng65GwI
8Cu2iKtDULvnlq/OSyfS4OvwgXM3waFxbT1RmvhJTcBRE8+ucmy0GUJVqwPB/9yGaSx3SUeGxUHK
rcpgsb98K+i22NZDNnrIk7A5OArpX0LpX3+QzrBTkAbjAb3MXTefuFBPPRT6N+vAFPmhuQjUTsTQ
fBfIbdquo05dVoujOScIligTO5wWwZe/AYJOSO1RQ4r9DGLZDzstJrBEONaRIy4O5br1Kg5ecB/8
piHFxoSkEiCxJJE5/ep2XY9n3dSMf6tOUZtbB2GI8blktiiL6f36e4EXpMv0+RVlbPZsXVeEY4lb
Y8J1zOg0E3PMXnErkMKKjid73RcGasG9C1m6eap/fSZbAsoCFHOqy7d/3c1tpGAF8HDEQw3nDHSo
WnLDySINS0o7ouq05zsSSutHdVvvRFenEPl2+FsMkifVz11yWiuv/l8s431+7IEcHWjz+D1irOsC
5QE8qox3FZuZFdjlkLvESk5cffL2/i57haXaCDSZbSbyRLBmVaJrn7x5lMhlg3e0vBijiY5sVu/f
jOfdgMlJS5kGD6mIoiB+wmE4fXQWxoqL2EUB9afHE+C+1E8TXOPx0fj7Fm2bz18GskFLH+JlopGv
Hl4YV0ohBP6oX3y/WJE/mbCnpOkX5DdNxqfRxcc/DOXJc2YXIBcVVrjz18xYLbt3w9GTujfMuGhG
TXFA0MQJOgtNVs5TzZnmyYaAAPjCEwh9zESowODAmXZrjQO5m5UErxLbTzD/vfLH5zHhdBHoJgmj
/J1tsTVOgDRzT9O/jo6FeU/d9BahmZyLxLucAZ/EGWaLbZ4bB4o2U1ov7mXpKVH/CK1Bb/8IHz3a
QeWKHc3NmYvpbzhrzin8vtLqld77rcW2rf+dRDzik7wNbn8NWWR6Mhp9KmH6VtpcMuYE6Ik7NY7v
G9JT0ZvDJbugQbpRTCWrTReg+5LIbAc96bMFUvjidPeUVoGND3XCGz9nx45nQ4sx58irmpAES138
M3/ZH26I3oK6dk6SX0qQkNexb1aZtf8pRMbmaUUIoW7s3JIht2H3mFVN9a/yk/c8rJYIIOfcwsAy
wlL0CNE3NO0olpYhsz6Jo4etKiw+kECgwei34KzU7qBnTGrkVHGup6P6pVJJgVR9MBhSBOJXNvED
9beDjeJ7o6IICIvugsaBpbZPUpKB7PWsxa/2LDa6aMHwP37JlcsplLK3xFzAe+D/rOH8vNlDvAHt
hMguAecaofpBD1Nb0KFBqfOJ48SdOurA9jql0OJugU7Mdfspal4qA0wqxXHQldgcBcW9i2b64rbv
JgGMzCyLXUYqbRG18OyYP1PslFX1vTe/tBgErKye15VcxXO+YZ55ETj0ki8tBvuSxXfZEIOv0qeI
/QQxDaITGdQYf6/5EPGPn1jt+jALHxDeyOKWcpaEbyIn4LSaqMXuZjUjPhDl+PSTWK/+dgCyki+U
5sLm7Wj+hDtVzkZI0ClaJuaH9TQyf+qs3BdG8UpuLBEONgghOFCrAOoRqG1kHPlP1kxV9Dck26Tk
JyR2/wYEmFmsmGPw1Af8wxoGjqd40sHMHNPDTyDQIpKgqyA5M8rhgziM6TNUUdy+v5BBYdpIkqCB
JSpY0evwgfDx4Kjq486CMCPD2W0/y8N5mftwPhrTWTDwwcR4R7RvfFr3ppB9qgzzryWdO2285A5z
C4foYP1vZAt4Q0iEyHzx+4sBOWmyKkp0A+fXcjHOcuoIKbBFkBOHY66H1KiLr9vX/591Re/UVwop
E4i1lggwtaisk/wfOajD6AaKqRMu6ts4ud+umaB6o2PetQyn233mlWUrb5EBGzgpS8cc/LcKk1I0
njMMhi1JrrtUu7qShJqTDHZHUIMXhXDJKFHEwikoh9REjFuxVnemgJlNvtxMoMAUHzMzsVCydTuQ
2jA9p7BFAOXoLDuvjyZJRexynAUQpYUe1vRFShZgn5UAuBIH5wxYIY5bAo8EMbJOAEe0CSAkLVj3
uq0YKXa6qvI3HzIYtqQNoxhpayl7KmD+A0+WENdJHHLc/6a98P+4GQyTPVEVuJyxDtXD3JvaMeRl
cwT91MIF+DbzuFc2+4/QV0NcolUAAyqextlXNAkTtenVSStQzKmA2F9ZRevcnhYlXCStt0UnTZGI
+FNFJ+JOrrRh73R2uD17CWPUqy00ikh+W87JkPTShpyQfriTLv1bpknqFFHKWcYsof8GccTJE2CJ
n4fHnD+SLrEyuxX0/w4+eDrf5mgXCT6mFycn24j5GsNWsUj8jAnZKY+h8h74FJBTkluvIo+WhXez
HVQHwqq5RQ5s8Ic9mg2YweDCBxWqganDVoKbPF0dzxOayAkWH8aYSMudK4zyw5Zmwt2qdPGbcA1L
GpgLnt7j7ZibtjqKIGXEnlTZMSkpHIxWDTPxCTKtuJyaUReMZk6UnaiD0RrW3EGJRGrylPhPNetp
Ogpu7kqVrr+YlwChyc4UCgI3ZUybOuPaFHgvhGoSjuNnXvewbjHlse5xA9wu24Cd08ZAQP0pyfm/
La2rlQfJs1XsM+4V2GwKt1O1L2YSnjGP6BqQPd09THbOsBbUIgOmzMUlI8QLr/09QMERkI8IASzq
QouqhUsIYW+O+7Onqkv3JETigTqjrByzYYjbmz3iCUR+zS4khnxtjgUT6ZG+yPlxXYpvsg69Mmp4
K82c3YEdYDemkqyPMbBir7SMwjx23RJPCV2VwVR93+EbS0c7Yat2DttA2kTMkQgTltFC/q6QI9SK
0bq457BPnVyP4aQmo7i6JPmZEWdUSuzUVewNnUCVkmdm4ruPInQhwF50f5Zq3O3bRTzqigdsLw0F
E/ZoW6GFEflwrV28MGSGohAbm23o8Ld1u4bcBfJy28bOv14CaqIU7e0qmQAtti3blhW/Yqh8Snu6
nJp6Qm5vnJJNsNTEUXhUZUla4B6bqjAhoOM6cCZC/rbeAP6Mk7Yby/KPbLEHcqy2RSEAWVPg4nGu
qGq7rIW1ML8RMpSFmyMVrg+gBi+wNYWmynjObhKg/2sVpasl5GTzaalr/9CXSbI1b/rlD0btrjwj
1F7L6od7Twm0IvlnKHg6RIcfeC1N53d660jRGzurOnPV6yuhAhhKv+zCmE2woqFiHaY+/6v691xz
WoW5Qs4TOvAmk5TghGjztqJYbFKyHqbX4AiJ+xcrAD1OOgiG7Dsit8GbVjmNa6cMQig0Gr1zihX0
+/+/CpvR8In5bu2qCWfEhQLIlULQdlaM7UGkmdn7SuSemZiUJLGLyRls6Ll2aPtJSymfwRykl6oH
dC2wq4/JXLh3l2Utuoxd7yHpOuXoCgz0A4vaHImxTLwSLeati1FbTwKksEo7heRczvIo/MCSavWs
sG2ZvfpodX5qtZLK3aCH0/AH5AlGXy1MtASkuDCHCqBWAiRh+xJSlB08huHZVQDQbrccK9OM+VIu
jDIHSXCtmMIb26FloRT2Dzhc8LKt2B7sg5g/cfPtH1/4WWO+GFKJW/UKIcbyPgPL3lF3IADAeScl
wsjsQd+MtV9Su7gcNdfF2DwOdxrv0M3XCD7lnBxF+izSFcSTFBnxMk2Q42fzump6voCaFv0KePJC
fTYHvmcoYkbICD6DDvsSgqfWoZhEtXEtC/oY9lvc07Q+ElwHXQNxRBxW4qHY7t644ybQr2uWH/ot
x9NVjamJFHRQWIXxgiiyRjBhnHSthMzFhOcl/SJht+WEjMVFMpEAydzqtZJH0UCXbXcYCP/PXYl/
wHqJU03/EstlQZqwARpBJzC9ccBMLtXK+GHSLm/FDNF7WTer5H7w70+SdqrS5y+7MZaYQm9qapPr
8tazBxzy3w3IQOaPhzEt4/RI4Y3/aJOYoe1elciMgteXPguQWztGuJ4/iL9R/aDnU1TBWpAWvYpA
Y/wYv8BMQa8IkK9RkSuMPDnWwHEoVGIDrVAsv+xnawHK94pgnYBmumtIOxrIJmnWf/lJZW1WIjda
ALpmHf/xFo6ds6pDHZGcNxJ7DM43GPoaobYTKxQnB/KMLGdX9VcFWWgOJxp7x8Af0IS2jI8+rpW5
PyVS7itwItWEdujMfW6MTG7mCAzNgpwryTtvqYkeVUIDb4oKzEtsDv08pZfzRY2T2KJVsnMm1lPt
AhXvYBF8MnFLj8nWLKuHXWs5IC4fnsx/1UVNDtG6fBqoKLNw5E3WG4+U/8B00mCsJ9LjZgwq8Wjj
ZFLSGo1h2XhZnWHcTNYwPEEb3/xfT56KnzfZLi7RSTPDIq+hmAf2OGph2U0gKY0Yugyzs50g5rno
EsrqynPkOx6PVpOISWgxa8jxRK+iKsxCwlwZ7hiMM28oKv5He0oLFT3mCt0mnkyXLWbOhUIfcXvt
0gd/KenfEq+dczvbbOuU1fFgdWlLXwZkc40ignpi/6DXmjbSrUQQMU8ZIVAtAycCXEnfJk9wvcq4
XeGNm6kV7OyWG4pkFipR7/0VPU2zeFC0+sHi5yb/na7qg46dBdVVPP9zh+CC4gDhCtkXQQRfVIrx
LBQHjve6EJrrvCY8paarOoyI+Xw+gFBSvZfPudLW+uqQvQqVcP7OZo+ORFNd0UyzsMfLUP8/2sWD
PvBRCz55EHdfA4g5zjaz/Bys9PN2hRAmy/ySToqn5QUCNf7pdhF55p5GDjBinP8G7LIrddMTtL/u
/Y744elDF45poD8uwEUgpIQs6t0rC8XAoXv7jz9O3Od3ZJEpKQEe6hggXH6JRHFtSD3bPasem2BX
DNcR3PYW99/7NToJSSVW3H2pYziUspW9YUoB1cB9HH0FxPk8/a38c3xtR7Q63uGFaZFxKK7VmYW2
I3xvZgnXnBzl8C7O6iJsmb44x5VBO10vZpTsE92ighVDiTU0Y2NOd3wu2B9CQLUPeJU4inoyd1PH
DWADtzBBb3uhI/U0piygtiE7CLt/jOYaiwt7XzG9j0/A7U/Nsm+XvJFB+QxGE/WssbWzLTxTWsPQ
98+vg9iwknYSsO2SKcJfMKXRfD9TXIkrWHt5H+o2bP8FOp70QBeoErHUEkdDU47wyXPigzliQ8Tp
7cYVky59bRtvkXKyFs7nMYsvsQl8rbDSbyEECd9oiSIPmSUj0CeDltXliKmPN1TNo6E+LgMoKOt5
eJdezDViKgd9LD/ikgavfcS1kxw5g55pP+h23k0DNZdijWz70E99bRIMf79yIy30tkw6u9XbYdoB
NqQdNJl/fEZuddpQ7EYTibA/1dYNROUjresx0L/JX65UkYQTq5BhO5lLbDLbdmUYmhxXuXLlFMsF
eR/5YUM5PX6RDUFVY+lX4iG77AjspSFRMnJX6exCA6sfthPYinKJfJljGAOSqDCLeX7eyKBZ84NK
c09Bi/1g5gPpLMMVyzY9Z1Ep50M2laP7HG9rOVNi4vYKrv6ZoK6jQ9nBAlXpiKVM9SF7wyuzJHOL
+ld6BsxYNNVDmD9IZ1fs9EpptuPE3lgnm2MlESR+s/7M7xhNoTUfCmS2jMFpdhHctcPu4EJjrw4r
iwp4NW3nIN4UdnWd1PX6gQEkRzp2SAYA9JUdf7ABDmTy/ZGx5bNT+XD2q+tQbkAPBqhgigPNqw+F
X6THhoB9V1BjqTmjFsjr1amQ1yW/xlVPdEwGeWcawOu1GK0go65Fc62FwJXyFbxHKnm/4rmJluJG
5xjmiVwpka/aCP9aoEJ6h5zr3LfFlcfjURgAFpS6MSgKXXslr9H1x9VXXe1YaQGMCsMj5qH1qNuG
bJPFZu8d0k4CWxOiU0YzSTfyNRCy6pe4T+tIiYCUxLlzoHJDs2dn3yILdJh1enQKjFPYq+hMHbs8
iCXlW6zqekHIPsjVc38Tvbr8tBk0AZOOLGnghuhhB489NTefv1yI1UYJPePdmoT7tk38RxobMi4U
/8xGSW6IOEomylAT//VAHaXFDQvzaOi3CZ0LogQNNKcszY3rWOwv07th5kot0aMi6o1uOvzlhOwl
m+qIRsp0m7pTqmQzmKpygHF/cLloakE+3PiAJKd7rX+PbtZRXPgH2Oce6JPBhPxkjtu2IxCd18fo
tikFHmufNpeXzBxzA53lVxwrRWlewy+viChbLKdpCmWVVQ9/3DPETAMvdYcXPEjBGbhRmsx6oicK
A+H74CkUZVZozP4JTDtTJkgn2ClKN4E6h7uggL1VwcOc0UALsqTto3MI/b9PLafXFL8AgAn65d/U
5+xna8HEJrMXlq2SCXCDXHttMs68jVWBKJDFDHj/sCCdO1lgtxM+79P9eQFiNjcHAkJO0W4+26CM
phY+REXMtNsd3oNoFcnZz8iehbrJI0LYFydwERu48K58ezecxL982c1xkJefFTe4oVmd1Ag/dgCe
OqC9recpG4w+znvOW/KcMaqur3BllrKGzgq95eI11SggnfdSRTg6cpwev5hJ/Oqyjz2/HmL/rVoL
o73WW4l7DGBxH+leVwv2ZQ+idz5Hy6znCnMxfwRShptBYp9cawfsOu24PONozAzT6g7XZ7mvKkEJ
WJxvesEwUlmKZMnjUDx3NQ2xwoHBMo4nK50iLmWbFN+HTHYK8HGU7nB1v5KVya5MQjAbAtt/+Zru
qNdn1V0WulpramaWZU+qMqdB7hKaqbog2pfm2ljipCmuluWlkbwkdYGvERK8GZWCMDzi6SXa4Ql+
jpZpt4A1IXOfdBZdwsNQjJFEHU/fhBvL8NGx3Lkle4jIDOlDMASBiK+siEGWmmljHxiLyPaJrjyt
6J3pkCvB4+sfJJ6RXR+j9v7tikWdM6uWk/q3E5875JeWOxMePdXgToeU/A/NaLSVbPGWpD51vi2C
cx2OcWhSB9XmFRAD8Gb8LFN1yE/9Je4PYsKAUMbzrZ8VPH5yKucX5bX8ZvvY62PtuXjMV23fHgzA
ioWXvmduo8+dgU39Y3NOKlBQF8kP+v4eBr7yogQLOt987+OL7nCmABjJck3+ijNclZHslWfRVJRK
skW1Rub9T+VfRkok6Frn0DufoePm9e1pKNZquRwI7urEz6LkamuVzcpezU2JRpNFFMXnLBrRHJiB
1E2WDD5kys+tNwycFRnHZfG/K1FPubslKIbfopqgc/KFv4Qcqd6iUrgoIMuX1ZbW4V/OoI6RwFNa
HejoFTr92hdfGdp7yw7glBOWiN9cjXWPZm/JcKBINpNXv6dUmHgTrv2ZEfIZXCskkOsya3o36s0N
3yhrFgbF8zh3orwaFhCpHyydSpRN5MezsBlwKLezJpuZEylPeXhei/e4A7J9z+Y7tFH7GLWqJWuQ
U9zaDxN35X+DEn1cvNfVw5HzQEfjayrFW3WgH35P7PyWsW1LKnZeVNwdZ177nmBKH2WJcotRM3Di
KtEyewkxamr/zi+D6CfSmhJ4kJx/j7NxkhYgxFODzptcsUVDy6J2NrcCHmMoOmZ/yO9NLeTuf+hq
1b7+2QzTTSkxQN3ADrUl4eijK/mbf3iRyVAupxVCSAAseVsLhEBAbCB8KQPna11bexyAffILHje5
y7vejoBlKQASQuHDhGAJ8RkJl5xmFXJiM89qltaoXZWGGMb5vZEweqfHbQ6eE7V/eRuPiBVCSnEr
GPGvIHSyjauAGILhuy6L1tzfsjweac4uLpzvo6r36bjRnhUBoj11hFZm5LSqAAoi1yp6qZxDR3Cx
hf2lG2aTECWzp1g7hREW0qk7pmO6LO+ReF60+PrUfbOsh6NCo7H1UR1SFmBGslI+m9fUqMOZQrSi
y/cv5GWUevF73/C9YyLZOyd/7SG5GbfoS0MqtHICyhjCyzi6hf7t1c76E8UVJSGnO/C4BaGgQYe1
bHejjTS02Jw32f1GU8Q+577C36OHIxK3zJG8aTCRsZR1b3R8z35Um+mMXGKYeEGweaarfm3nx6gJ
KD4W7UehUOAnKq+lXh6Dbz2CxC/I2Ekwk9amb1ZfmvaJoVi00PqmY6G3WGo4W5Ht47+LJGkYyv+Z
o8lt8xjNPHcOwvezar6CZCrKJ70O6cwTWQuKftarmpVTtH8e6tCwwL5sOhS/31h8uWFNAfbzMolV
3d3mQrJy8jVWTyn48UVUfNhe9krw1Em7vOoaurI6pyPwR/lWlKZqpXFPaJZT3JKzp6UiMo6IML/R
83W2fviuytMFLZff2dFx47NH6qbr1dmY1iXtDjqnGsnlu2S52+JAJXHiqiwP2Xv7lhcKzM/owZ/7
WlxVCghImRFcClbzyxpMUrfo2Sp/LFiL2d9vkvwIGV3fSaRS7qe/4/L8WhmHGnbXKujwk+YRhI4q
fRAY5gSrevM2D/Hd7VHD/B54xZJ0h693U7Wm8V4kMr/MrAONl+GcMOdJKX1BqbPv19UqsYljAuvR
4lbRp12B3otHHrJS2X62Yi2g45VrsG+ZbNBPoNTQ5kfqQkAbTIVrGPd4oL/ZFU0xAgZq1eFP2M+n
cGTYpQp70hb0tj15bar+5abmU7cQOen4zLjQBTjaNvwG0HKoQLfrisCOYzGaCjAjLSrO/Z+B2+I5
ODSYbxLF5Qqytalgvu6DuuFqhMpkAgzNIkKiM9XI1zOfmiLtp+Nimpjfyw169SASTcz7EZ10xHIP
rzD/oOf39i/IsUSVu+dZ3HSG70P9V5WhKDcxIwhPpKGDPy5r7GW4XJ7KcgrV6+/nZSrNsixRR+bs
7ZxVu+LdrGhL93vfTdtfdA3CTD0cQi7VQIko9Hc4yEoMpEVRd7iv77g4nK0qDWslSsYt1eWAY0ir
WGHO7vMjywm+HTETwAijGvI3W+4uqdLmsFSlibei014BXCLx6h9DAl2u2zmytnj8LL+lmd8x0xQE
ENKtQiL2feNMKaFgfj5Bdi9K9oJPKURY+Q/1hK7kof8lG7olZn+cK+nEd4+PepDFcO9OBXvw+bV3
vKkujbakLJHi1SzS6DKTYAxIGGdOayvdBwwj49s088Zne7eQ3ZhpTZLLG3WMsbfckjFaN825VA6c
u9sK7AyMN0zyo74fUC1GAAdDDSIpfYKq3E/GKvt17WBhFNyBAQWRZ31XgfaSHg6VgX4XtGf2Tx91
oIhbRRRd4b8kwxiAyMtK5959QDmT08x+ALIsYrcWyvpQx0AY90Wf0X+dmqUAWz8H9QhJVFWwFLdx
RJ5xIRPuY31EohR7Mo7a/3U5CbISavcxEao2Z0qZ74Ph3u4eUQFXTAVApCPOpnE6kOGeDBymGh8b
eVew3HL+pglc4R/d3zltZWeARkDEApc/72WKi1V/3rpnqDMZdzJW6d1ov1xvVX9fIumRHJ0RPTpt
W3+9O4p2PAek/lwmsGu92Q5zqr6+lww1d/qYyOME5acV0TMsZ7cpXHvXqIKUqzn8BG84pEDr8QlJ
QxCYs0PkP5ydH7jO4OBSLZ6lGD4a2BLPSTnG7lFhxH/HexPaq+PetOh/dxABwVxE5A6vYL1Rc0+p
T4WXS6oRuShHs+SJTom04cUAas1mvHIGvmrn3odKYs06ZVpqxyqWlBHlrcjiwkCAz9rOISfTvrGK
rnfy5rdqBQxhRzZ1AjnMHLb5FAuMxJBsFQqfkwJH6vF+yP4oXDAs3TaZc4JlzwIQft1fL7rNFVl0
6cQG05YQs6U0ZdACNrqfd33254Pl/RXOaeh487G3Tdf0UXTTq/B6CtPJ+fLDfn7a7wGuV8z+5GDW
8dzD5Ig3simRexiIEKxt/wijfkXN9MSvc1/e9ILaHeNmswR+okjO9LE8WF7dZfbJ0Y8lf3ZWyqHB
+VHe3RmhCqM0IsiTcjiB7fbpH27zjo6F1GhO4eluJXBEmDhV1BFRXrBHvYKGRtLbm4myeJ5aQ0YD
42Koj9tgTtKrVj+V45cmlpfrsCQho3iGVd5FfdnKVbf/JLO0p82xdEVMOkihQwH6JYWKzGi3kOMk
m89EbQq+YPY0NZ5Jeb9EkwDd6WWCrir5SOT6fbUEx0syI7oFogaOG4fsOFoWIEnVQOiA7sNTTe9M
A/dtEFoqpIjtEZqP/1Chnauf0SUQD6iUcEmP9ObrnvwhU31GpGUuIkljN2kP+5z/UAY9jTNPf0VD
C0j70HqAw4L3vazGtfQWd0/4D+Uaze1qFBgn9F5KjkSYWMv42IR9U0GkIfTTuStf7/9+BuPlzPmg
MjIwjwgz9qThkszh6hbJpToTXaB5zO9pq23glLbmWFcpdbEpAdl78V6J66soQGRaB3RC/q5kaxNh
Hvb+aJ2vL0O/yB6KdbNV8ZWGlV3jn3Ao46ULyKmXvMFwIWp81+jV1rdrFB9AtUiZ0/Da7cu5JxVs
NGeI6wpcZUM+AxptxMDKHCNySU9B44SkmrsxD1CJqMMM8UCtkdMhXXNQH4ibNrorFJxdXbyhEW+1
9pmGnL/ho6HSdiaamjYJbGfIgzlN465aGB15eoayziLJSlA1abjrQkd0RJcsaZAoZf2GKB49ZmQp
50v2EkdRqDCxZsPLZrZhsuf7TE4/f2I2tIi0qEx/ByZhS6vr7cl+ES5dqIMRWCVAzAT8SJJ5QQ2a
fwr+J6cUqPV9bOZ9EEulBHlo7AQcddQeGzGswUK8PtCQgl34iQqhbSMb+fYgyiU5MRNJUNGrB2BI
vZroDiVZTE7Kz9vpbwllCX9kkeJR5SUZ83G5oFzXrMNJDq2oqNtPqcLE/K5ebs9XbZ95g4uY0DPs
fXZmXL9m5WK0oaJoLZoJZTZ07yIroECQd5eIWNbuiIw9fiZkiefkopKde7YpegRh8OjsmSMoM4uY
D9yTNYENgsHZ54bhYcPxAt39yXtLuIL83uOaWoBEl+A6ev7CBXmocF7GIqX71kiczoM4NA74rc2w
iWhHkcvgOb4dBA0HHJcywM1G2tT93jPNur/zm17XGHC8D+p6yWQBqPCETYV5sgNe9sSpbs5UIk58
tfWfAeybqQMG9wjMTUN368D+3GNEG6xK4gEvpfg2kR/4BJd0UHbT3yiLFzNaHQRMIDnxhJwgvCwG
iGBkR0U8CX6ApjSIlomRXXI2phvLvH7MwOb/HHO4FdscYFvn1X9vvOc0+oVeWXdgoL/1hOVLGon6
VKlq2OQ9zgf/ZKkFiKoOw5ol9wrMiLvixqr/UhRBWrP3LCvFTdSbFJNavIqC59jYAZgUW4rxrMsa
i0XCGYtEhUuIQGQoUJ3UtIYyxyOAzc6gsm4vGMIAF/72wKwTPehtodTCPovhAHgsHexSlOdetLuL
VNGo5UEis8iPCRPKq/8ZZ2k/4CyoKQfIzzEqChUotFuCx9w92PSr/L+rW8SxO33kBmIwg9EyvYTC
tB9knLpVQ1st/6FKgIJdP8jy6uA1qdMySqBj08Olil85tmJw2YfN0Xbnilqx78tSHLT4fZCiPbFp
QLBBB0TajZAh+T6TNed1Fdx1V83SDmKUAntelEpA7UUdtLrmt1d+IZybcCXsjq+4nx/KkX+Aj1CQ
vhbxKHrspk2s5f3bJP8EwuUpPzVIjz7WYY6ljhpf31p0kPmh2dTgJvYVWOSPp8R50WluNgSVh5w0
r+M/LHSnl9yU23IpU3MOZ2gEtjD7NhSTjcbz3AdN7HFtsc9vhwPN7h5eB441pQfHtVhUywn76gp/
fpwe7Me9kG6WyxUkSNbhyQGTG+XKf81u9ymSu38f009XQQfje4Dr4qcRT1vFVHuAY0uOyStpAIeG
14N2e+uVfVZK81+nK+KfKGo58dF606zvK84djHSjBBOvcdJmVeXnRIqcLs4eIoDh88E+461mRo1h
sJhsejaSXMzAGJkAhk/3nR8y/X6Jr4lZr7drWnjb/F/nwVUOd5q54vYtR9S4BgLe4Pp9ad3G8ilh
eRKfNEqCgbUT1Bp9g5qO6rVel8C966C4Nq3b/PNpdmH215KWwoVW/cF3k2P/Gv9Zdm9HtIM0lUde
JLeGgxQQhXJqumuw2reKi/WStQ5fpni8nmYJ/H2X0rBbToLnj9c2DMwcDQJbqIEi/SUroUDbU2O1
fqU+i7i82quPRq0UvjiB6aneDQrmM/93964D/WzsGfWaELz3j7Eul+lNsUSN0abfSSDvPO97eOzY
tw/A1APRyBC1pYmViMxh1+x0Hyyn11umqVa0GIy14rBxTLgGvSwHrJFBqGIxbh8FrflSrUM8q2if
qNrKFmlrtCwCCGuaHucvBsg7Pe/4XxYiXA75FRAjFPumIjJYsIR6B9fVJnu79yn+Y+9585MUXxdU
L7GXqR1LOmjYh/IaIRZ1bkOFacT8AWuPGFnNTSIgz1DlojZHm0Dwku8JyFo3gPJxPR/lglkYoFIe
ld8kEO8ufwq1KMitgG6xNygbK/ArkpMRFvjFO+CrN8GybH1eyORNHKP+eXkxDxVRDemv32jcu8vx
YWFeKDWaNN8NE+5Da26Jrk0qQxZoIVyFn/+JN46TuaJ76Jvfu1OV7I3HwPNRmQHy4fUO+Nrwz3SH
KhmkMAIuhpaeRAl8zR0FOyyqy8//RbbEX0Ztbzlw6jVLIFu6RWs8bRvAcetnYYr7ykf8tIxglLem
C9nY+gd0n6FpkpNcNkC5cHWbFuUqHc181B/GvaR++mCX1pkj0qJ0neoVvm8haozSkaO1jDEYlYTk
/Vq+DOn3CaUNWaVJAAipoid0aTpu1j2CVybhmAen2kgG6LTZzl9DurkeDy79cG8FLxwnW5xzZKBU
bxEX+y6pedtvwA0/yIzyPg+pdf0Rea8QROEojoT3uNZ63SO7R8lZ3wnrWwcmVHN5byfygEPTgvpX
b59qsC5fwiBBzPLkKFd8/iZkYcXOwAJ8anO7TgeCQQ3FFJnHNqN4cOt2nAJFCkexjfPqDXON8qm5
JVGVevowb5jFaWUeVPkV1+rjNuPNj3asH+ehIZS235VE+3dN+syPE6BjY3CbrMVPBQaXQuPC6j4I
+tbkvkEdZriy6MX+boJA7GbnAe+YzrKOPelpbmvN+gL/KBXl4hUOjVs1GwHlvBMiiCbmyX5nPpz8
159rDt8ebAWuN1kla3mVRDBBL/4bkiS120r9ulVkEU+0DBzkPPg1zUARx7AGS5MJQYjaU0CqKsUD
WKcPKBqzFXPnlQo4dij8Mt2ZlC3xM+kEtim2vCEYDP1cPcpjXw3oWMtC+S7lMLTzLaZHhz08vXhD
m8Qg+Dj57c43V+uRL132ey/d3gqGiZ+RLAClSVCTKtm24R70Jh7R5f6V9RvN3bNw8DKRoOCQtimX
1fmWh6P14HhuYUMR+k0ZX1nme/Bs5bHHF7ROYo5vuOA5NbSLaDQj994bv1gmIZonFwP81QWB6E6D
12EGldjkWDuPX5cK6lZrB6+BWlidQeg+x11zH7qDvYfSmlLNF9GAQxR5lDUQK7b+alvckj4Rjp+t
wA6bcRp2iYbr09H2uKF0hoEJyTwVfw0QvyNMYhR40BXjltRyJDOWP6kqVv7IUNdHhJiBBOmaCjf5
Blray8u5DZEVwMbiuKN03FxxFsFvj3zqij+cgq1863joaOIwqLDmfRywKQ6dvirKKVy/eutFhj2p
56R2clot0BU/nN2/NXOnM/DvM1mk4hwqGlNmhjn/BlP8Cu4RYfTyVWx6dozgcAp7HGvHJu2QY/zi
rF15ZcomsLjpGww+H0MKwjnqF20MvBVsmO7fwY4OHXM5pWC0Xohtr5GjJ6SKWAEr/qjGJfQFKW4E
nFO3QVlFHXNKNXAYohAwwZczrdg80tTg1GwKdu9r7JoUHON6ZSTp4qWmPeExuf305JLgAK+vUcI2
VwtN1Miz7LHHGbjKNQDZ5f4HYkSlNPzOPcRtA536jQiKssliaZ1aP/rxAWxkrLR7G2g/wQgCUK3Q
ryEUmWf794dMSTuafDrM4A/pRgRYNUOAmaHD4rK7X4RGxEL3graIu7ogiW6x6Uvf0Er6PVl2Asbm
RQfXkMl8uV/L4Jvl7lZGKRMnuJ2BoS92necKMfVk/DWJiDanA2fIDP1VKoxK0NAVBfu9yBQe8WBB
4a1TYYNcjJEFGo9wBb8we1Ss/Y5cy2XlwrAo7T2ULmjlUTWSKHb4qHAAtq/v1aTEQLLbYXft3Er/
Y4Zqg/T3a/icSpxlGxwFA4FHkjZafKvbvVVTHieB8iUXkSHcT1gp9rkY0QB7E74pLQmbe+Q7b495
szfwDz/yHttZ3hZfyprOi5bTJvvkXUkjmIht7tEYUCYUHLDQmZqVW6nnZRb5zGb0NsAG1SwTAlLb
gojHQbNMKsPmLm+4DV8xqtMxxp90r5itOWq0miu9U006iaWHIFhMAjz4SO7J5bpCOCF+1gw4ROXG
gxSX5cRbsMQesFQzLo4lIBdGqBcnLItTn/1PicM1Rf2ARPXAHW2st7RK6lwMvyDLBY0CVRLSmroZ
qpNxmZEAzhZULDltsA94sSNahyY3L4UjKCsQAPHqNC4XlZia5JUe9QpXL9wdQ2Op9GwXuC5WgvPF
NLC8yAhKQfFprNLwQFr0YJyxKRaKcWMKeiHyuiytsF+0At2S6Lh4flSSEIRuoBmQPsPQrVDv7oJa
w2tGiyskNNSPe852HhT9DZHfFERuFPyg00/KIWeSdFSd/yS4m9eaNZbtvkD4S65PI9qXsShOJhg4
lnPDKqFC+3isKnge/7nGW2HztVqsq+CSMRuOGlJSdZIdNyBvum9Jt35+m0dFPuMpIgSFh+NwfHx5
jRcOxaYeyxDoJTdj1DLyi5x4QYz1qOvh3q1FKW8G0kKdv+qhVyG9M7lqmwcNYJ6xyxQqmxIZF31F
gATlB2sJQlchDoEpGVW+ERI06YaAN836/wc62pyXkgTXeAkyvOq/XY8tEhVDTT57IQoJbvnDILk3
Q3DF/iR5WOqu4eLUiP/r61wD1LTZKPkQ24lP33qlq0RDLvCO0AZSgbbU2dGozTNpvo+oDixBO1BE
Cg1w+YefzptnX1zGo+9BYY/80PHucNBtHc79FLnfKZK43APYfb9KmBuN0nXC3LLFNMmTL7tXXzEE
t3M6MOACQOxv4wt61371OP82padofJgHNh1BKX0f3n1ltfPyyasj0tqHUgnq0S/kjLhHlRLYXtFO
UD2ndlzQsmHOpq5RqD4KsISACbVg+drMPGFEbNnIHwutZ7fkTfGWY/opUV/cYjiNx3NsWT0zDxKz
yMAhu3gW6lzXw+SZSTkIVQVoYoaqQBUDVfOTEq0SI44eGKTc5KiehAcs/t9plp2pWuHqwV5FIxhz
2OgKVaRFNAdodWD5uXqjCys+t9dFX2VDUX40U5bVEvqmlWXyPVpEunZNUwNR5x9vpi9rN3LMr8t3
jullpChgvEK0pWibgM/3jlYHK0FTYa1HFkIWP/N4V9dfgdF/EybrMQlOJWJrskGHZaNMvVPoaNQ7
gAcq9WOxcX5InBfvb0+kwpIgEb1mUYfDubqwcSUWpNpVf8tdYPfSB469qt9zrFZhbd+sMmBa65VH
15Fg0MWf7LW7dZxyCHUeKngclPG84nNQR9aX7QKVI+kh7tHa+nuukMax3rZNpLd4/HdPRoeuIa7q
7jmfV89R/h3X4hirqmUrRgni7oAeEY2f1kXjWAHL72BpHAsObrjiz2QBFDPqPmSE7IK7ndKf2C9D
o1m+GHqmdDuF1Eb4x2hcOSdaCJnY4LLTzNMKrvTrZAcCwVDKL+2TrYssxjFJ7dkxqS3ENaJz8Cv/
uOBBMajmNcowFMdv+ZKyXBSMHf4qiLMGyaNMYp0vZko9Rk01UM6Qi9TsQqfFAL3pLS86azIgGjFM
F2UVVKGR4NPkgB218iaiRw0/zRUaEfIDtvZ8e+vknjvBrCVEAOsL69YpuB9vxdGBQuEnRrXFEap2
H1cSYU8CklQR3tnv+jO0fF8GBdgZnGZkeAbitz9SA2ppcaw3+7Qbg8ZJeUn6vZd+owk55QBcZWna
aKZ4YGzsHxOlU7Vj4zz77zgM6w1XDzJxxznBpT7hJ4eGDorEQf5wf9f3/uKiGcOwzpEiwPhv9Wdn
dHU3REYvoSln5CCX4BajrgfRVyPu6DheES7c/V532Xq0u9nXlR0C89RjtQTqvGhEdrlwNu6oO99Q
OqJ4XgC+zIyDF0Q/1qIkObMgbLhkihVTKEBSAseeJwH/L/7bny32345fRin5n+VmQY+IoZBBR99d
4/mkMUP48y7/MzJ/qyMlLDWmAfV6FWOrk6AeM5OWtGKceSxfZIPYMLvs6d30zdD2pbih4LqjukzY
kA9zq0P2vDFU4nc44Yjsf6i5pFa9RW7yrukz+ZgcvvY54a4NSnnm4j4ThIh0I16OxDDBUwt8d1AI
CYH+9tJb0/ea7bCz+K60G16OfOJHddW1O/JiaD3qUN7+LAG+VWP8UmC+27eYUJXB7OXuYoaBhFtc
wPz1fuvB1M8+FHs6q/0KfYLV5j/fXJzmYT+cCgdkf+A/r70p5Vx/UuiAxDT97GFnKuxxTDF2bSbJ
TmwJUe+Zn5sy84APcx0X6Ww1VsG2/1iM0A7Wqx4jpKUl2cZDRonXoBx/m2//gchKTdCa+g7OlHoG
PcDxT6bNLI2rSMglVg2k5OlN90CHMOYcQPvM7nyo7hvt6DVPQnSs7C/pFDE/KnFPoHWuh9a2BBJ6
2yjf9bw7hac9d9lpAsOcNzLoko6oXNojNBGlTTbzo74s/yVaFMdzHlqPJ1194YT+mkiloJngWTDE
U9pO3KxSkQQbHbPXlG5egIJ2S+xmTgD7C6y6VCYM0b+L+YMIXwzvX20E1nWQpvVDcHmaYnTVyGte
S/TtrZrdh0Mdw6bl0Ocgfoos1t2K2l1LVVXrwFGLBpupeeKqjaQ5e9Opc/V3qVc55hSXtlxekG0k
RhnmswdhLGWhBrGGG+6XT+rC9z2861IN8jpGKi/qtxw0DyyG4ZUPYmf4flE/koVDSOnLftj/oyjH
n0NCFqJIwEzZaxM5qrsB5b+zlMHHMeuzMqbR35Az7Nevkrzq7HGg8KMynKFYayH/XN+2r2hSHDWv
kE4DqIWjUmn3G/HHUf+1I3dRsEH9OkurxTe7u6ELpilYzc5eQ5+0G7y8z2HTpQDXhGz2aFRVXFpF
IbiHuB9wfr3hS8OGzBpz33pZCTgMXTwwajmwwrd66j7I9pkSeErFqYoKpS0JccRfjwXedLjRpRRy
ZpDc3CumJ0tTJQvnUvD2G875QNHqxQWG4cYMskiBIjQCtvrvUqE0x2lzUyqA6CQajTm2GF/QbGBM
RKAT2I8TxZQ3uwaGt1k+dHEFIuUY1pV+bBGcskzd0eivjhTnqPmd6CwnerUFnXURy4h7Dl+9hpFP
yJ4pTWISHhA5NCEPaQi4VLRhNsnqJlY0A2pvo8/P6lf3irfscouWFYmw0rgEL/ZG6RN6R7vAfzo4
rniyyWymqZn0pMSLfF4hBEORb86WVDkxir68Aejifj2yQbbwyEzqINgRt0flHOvaTxd7XtGnO2UP
ZuyBWZM/II8J8piLCGxgWFXJWbb+qifOILTet3GHzBZIofDke4r6dm3uE/HgGZOwvaW7z3i4b9+H
VZPgP19oZWusHci8oL3q3HW144tibiCsv+2FE5wGCb1vkoQEbVkf/lyWEChRFlp+TP8NB7PsJdBl
ObArLj0a0FXXQvdFcWKo8uxi+Op0u6K9YqBjZ9rbQupLpefFxhvrS7tsOY37gDe09nqji3kZrxY7
un6CB9htLxWjzsSsO1luM7byrSrNsoCro09fM05gHAE+OzsQPCntNf9shejh4DiJ+7HllPf9+ml6
lItXB6svsiW4AdMWlW4eGF1q4rZOWzie+6Jm6vq00YCB8p/PnrsgmhXt27Zm0KCr2mbzmmaNZWeg
PHl6d4VgTKZKUHVHCwZ9VQZpkYYK+Z+hSgNXiI9dV/EzKM86oGucZYYjNgITRDUdcAkkfbTTY15n
GGGIsNtCCDrZiXWXrW9MoAxuXabSnI64uxNH3JeLXuTZFeVQ7xvZARJa2VMJWKC31bOXS//ZtXep
QtJa5dNYs9I0dw20Px4tdjYg875pyQrReXSR+ynKNTHydx7mpLhj35ztLdD/onijgO/Bsgut1M8F
2SBDA+tr19m3pB26dMrNW7tYWXg4JBjW+94yD3k5dmyXWQx7aI/fWw69yhw/XOcGogyPCvGLZvlp
gN2Jz0NMmT6T+3VubNNiFdro1tOd6zhd4o3cdPlxAgRXoLl9p/jiyWBJj2Ll19J4SD8Z/s/xbFGV
TVig378zWSt2sy/Jzick1PcckTGMmczCCvwEN36tIcegaZjZd4/FxeV+DYLXIVo58+7PwgX3sjDZ
pNMlktrRAoOFb6TUSTC3kR8wx68K7Ajms3bSJK3STgDusInveFruIJc59gTiNCcw4pMsRp+peMIP
FNdWp4RtpYjGRdsWEoktc4mL4PPJg11Xf23okdye4vmH74IyIq1mvZYkKKdHnnM1ko5oFODf3gqi
rPiW4HdK3DpnU3VLB0IKhy84UCVmOCMqev7eOVVUcazv37kDWDvHtDaJz0SZSq/xv3vbasuh8RS7
Z+IKxoqqZmMaokaS7sBQKwH1X6ACKokSu8+w3J4TOaKdCNPM1Ask8+P1crVj2pQ/yGJsSx4aDV/7
6oJJQ+QMQnhRefqZcE0f5PpLi67rcKTuxOVakujQ+dfK1NPonu8JwURax9HbITV6iAIYvY9I8eGA
J/txikJ2ic/+BcTHGCrUsoHvb6RtuSog6cNkMsPV85q98v8OPAB+9nHk1L1hpnIUFY7iGAzWgsrm
j933q8b4WP0eYtpglvPVGwH2uqQ+SZqB6R7WND4UZwxGT825v6w69cvjtd3GC50QFIeyOYltMsiQ
fzgXqy8iN6IDMKKZfHD+zWmnmytQJ/TC3BsMYoKax6ZDQU4iDK0l4zxJLLcrgIEXMPvw3pBV3lkN
RqF2E92HDvarK2AoRU/vUZ7PAcLUPy5noDLfRXxIEdYnZTYqoam/18xgNEXa419TpKSCzY8pXP7p
ViHigDpMQpOBMa2W7wtQle0Mt/9soQXqcQJ0g4+neW/vSK7m/TN6wc5d+nweEX6rxzYtSEH2Sycm
g2Hf+VTYP/w2Yc6AnB7GPLfMvxBXoQE2b3cWJ/13FFVsECCF3p+zaijosF/wK6I7jctK+Lasblm4
htEc46CHucwf2klZoeCJgalc14wKuMrIGVHupBi9Rl1KeIuiZZD8boY5ct28dsNKQSP+cojE52+k
+eiHp25uVbMbQnMnPAPHUbMemOH15dGbC/zCH+gcGUUfdFXLoU6ctDNiWs9Fh9NgjmbUf5ErJvtp
57BcdO9MIibbwizo/3g97xBkSFyNsM4NTX3WWGQWvI/QBPmjIyohxmJ9OjCUsS/ROvpkPdx95FIA
n/3shTmnfaQpl5QuvjTruIZ0euX4V8NqHOo1QBOZTRj0gJo5LrE2kXhNy0S26jm6taQzzAPfcYWM
M0OnSermtAP29xDGb/knGjP05tX2JuJyjbbRF4xv+vMiGBiq02ZHEz/s83DMObyBhN45TIPCcC+m
jRaEOihkVZjXwscuOco36Y2eRgeAgkUqwDxf8ocwEkR0LufoshBA2deQu9PQqUq9hKGRR3x/GepB
Spuf7MN+ivmh0SlIJfOmrg2+iPsjamtQ+GgJeiuyTiaeBr+xvPhOGBuzIgn7omo9xXMn6RM2WihI
2WjCIsunXiolxxQhZeLcMXthaOubYBGDbY6DZTNzWeD+DuhgMPGbcI5Fbhk73d7tUNQwdjE8tBPf
vs3NynLRExpi3ye3xkC271C6GsgbFMNWEDo4HADw4hbi5+eMbEfkTQJiqSiIRoVvuHMB6p4EOfsQ
PxCMk0guKvFqfZnwUA60HSRMIrf20rRCV0PO3XmL1ETIxi3pGcqOquLxPkmQ/dP99KPANY1e39qc
pNW7BT8nJUW8e1Q65G31U4p8BcxKjMCXEsx5jiGIM+JMbomjfZM6iP2YiqNNN610BzYDlONBeRNT
fFVQcvsj9O5gxWFaBDm+RD773h0Cm5RzsJVFlG3cGGwZTnGZqDA5CMnItdYPHKTXwOb2p3Kf1IFp
2ocpb2T3IJd9mw9RpLROLSOMSoaexUoblGfpGbCORUX2r/azqEVcOu465u9sXuZlRA95JDuMFH+e
RUDVsGjO7bkjeIzHOZGQdoARwRIW2thn0HZb9oNSf5BwhghFJu1qTMs5bsevjNBM8W2PcgGPKOTz
IxNMUzhjvHQjdLtmwrqqM7a3tf5qrSTFQinZLzwYmUg7I5ieiN123Q4Ek0hpX+wz1siBzceAFK/L
nTQTckBALoLERM0u709ti2ZKT7sFX/HyWWh/C4y9Z43V1q5rwL97g1ua2lxCAwhmFXJrI0BM/X39
WRabPsXlR+ALvx/KMS1v+yH1i9vqRtj7Kov3OqlzMPDBHLXFYk1fqdYhPY9ncwnni2C9xU/btO1R
9ZfhWYB6cCw6DRNqhhWumLs79o9KfCrGdAND6i228UHXjzEYMm6X/oxtWHVPdp1LexWYcuEnvZpW
OQ/QBjTRULBGdwiNtdd7RKupaT76wT/4mP06xrw5mcYsbu0QHqywnjCiOGwj+0JFfHaawBRpZd+U
HKP8IrwAzh32H+3VarK+fJydV+lWuhUgUTpwFfniGvG0g2gF24GCrRxdWOcu7qGmTlb+P82qdvQD
z2lbqUsnyQWyloxBenbr4A2YaERL8NMKpuL1JqogI/k9zu6UTS4Vdzvs/IDdv1hFmMUVZhWb1sOO
/4TlHoGzfMjp+wlvRxyMxAWM8sQOf6aEWOCxjyvH7fMSBYVntaid/CtxJYl/hV/VVkl9gI5xcVjq
OEtUZUeaBnh6gtokkXmady/GrS22mlBUPF+SWuOB/XgQ5PqQBmQmJxXAuJqSIT66/DgEhykCwOS6
caSeHv6T46WvWVsQjTxnyILn1fR03jE9l10+mnUrhGnGNO9unjk5R7aXVXKWUvm51LTBDm3Ccitw
58laQnQZgwQ46nv5FYITrqZ3KZSDHTXlrFdsYR9ziops7UosZ5LOXxf8l2GTtodZdR9atR6qXzC+
OjDx6FReYykkYJQ1MvV2PuGVTf+URpDfHCKHTn6wqOu2xDl2PQ3y8in5+0ApG4K8ZBOgCdEJVMyI
qqkA2S2HEYLi6jMrm603MIfolslfbolZxwhQJX3fRX/hTiMtG6DpJ6aMmIAEM9IqBHPD7TprDz3q
02cic0T++8HbFmT74DGp6RyNdmIMibDmb5n3GdPeZ5FlYH18i+pzmLt2teInBtRxIkFNp+dh039b
JE4vplvpLZ2svzWxf/s+wd5dQ3N5inpqLpSWEY7fuGwBmXy7zx+OcfINGjdOuWrvkiTwPq8Owxiu
RlF459qIhzfrxmutlIMnsI18R17Wrfocx3xBdvmEB+xwoEmSrO2mWzWQ8aC2Lb/BvTTLJ+3TkCxc
5NEo8jsmYP9OECWLtvnl7lcrJPp0uaxynVb00/VFNYhUJidtoNXDiJ99COWYdFWHjAOJGjCzBk4Q
EN77mXUoMWplHtQ4Ka/cXkHg0jrFVYoKoBaRiWZdxljLNag6zaSGtfb0qINcNDmaC7662q313Q/k
VLjUgLuWMAxsUxsKKY57Dk57S4eYbtLthId4K3IZNCqq7kiothwzn7YYdoNHqLZXcroJm/b8V/AU
pURxyo6Qb1vHFzTX593mmaE8AP0Upw3SluzInQ1RkWm2xXe5z+xbRVmYGbJzkkOphmIpMI6H6thR
5crFOUgoVB2t9zTQKje4YNZalP+YU2js76jabFor+erdmxzbfmkPDtmz/8gd3H9pz078HPG0h5QF
R/BYBN2BuRb3LQ84vriR1Ly34KAZ1Te+4rPbR2o8nlCpnYO2WY+Vy0n7oX6uVpGyt7lu/SLgGmm1
EgkBHAQZ/tzUz7Bgk/eLVuscOmnF3MgzSJ4XsHkZCh2Oyq4oGhQY7nZ0bVqHjo8KmFAHUa3DfYqC
jC3ZjRzp60pBkKD9eJROBZdbKF72IeEztZxfmFiagD/QEYyVJhoMszDTHhCGakzGnX0LKDFnbHxR
so3GjDY7vhxIYBh5glnWHLDdp0bErN76mXn7i+mse3XTbq5L8sEaRnG+rRmoSNarE2aWc+DBAw++
/oxwWGZcazHdNdfiEdHfvVYQ3Jke9UPKb1rWWrFNlNrIkiSHnsh3z3kT3QdNQ2aP0vPInsW8Dm+t
RGSOiZkyby3ybUoRLi9tOzRKCLbOe8fRant0gjmXk4/3rzxBJWU6g8L2Ve2iScFeitA6atZWTXPQ
aJHoXFyGJ3tLe8L4VYTeCDsAMckhNHZtFQTO6CUKQ5lVvMkzOv0foBluOP3zrBaaBXv47yX0o0fs
e9QNDxdwqARc3/HHkLuLJMDaVpAl75DgAGRCdSVnGDjLfQCvOjSMGb0hjz2ENUpW+fmlPTdq7J5d
S18A4kGbxFGSvggfZQ6xG3OTtos2iAerbFFAiJdQCPNO+pHOcJ7rylRpt4kcmFv0fa4nj8BBKKbI
FhrkJb5IsF5R3Hs7dasfgCmsgP9bz5mjlpebsyUwtaMe+B8ZAAgcfG2M+IzMH256qtBpOYfMDP5F
3QjBpLXwDVX10PT9O8KV5/RiYATFxlhxX2LyLmpIaGANCLJmTHihh/gc4Z1ry/OOgkeWabbJZIhO
Vqx44nalNye40da0ykuqVH0Vbnz7NhVT4YSZgHUc7fbb1M4xrvywDbp+1k8nhUmhVgf2cRFbQa19
KKah6oUFmuJvV/NKXvHM5ASDfSTwc7T0kEwtX7VUx/vZ6/IopUgJqL1fcPHcn1vMRysv63h9l8Hg
dxRdq0EPqbkD72fidT/NZY98jagN0ClQX473SywjKWfjIsfT7QYDkyQdti/3VZ4zWDx2WGrovUan
6H+WG/cNhYJVtZ+opL2hQTYCAxz7TUpZgWTTASx06sEkp8vd/ZDuuQ4bF9eXpBhmQERn8dfWRNdt
rnhS5NEQ75PBSKZdMaK/dk0cif2ykW0gefnDzjfhKyx8ho4cOdsYtIDXfCpuavAyY/QEWZOWZ5Nm
9H3Jou3H2fhy29mCJc+0v7UuWmzWQNPeCTJLnFsep+8fGKRRXoeyj0m42WkTv/7RBXGtKgmrTA2N
/HMBjEyC3re1tnyOieacN42yjrvgw9gbEYP/gorZxw9IIHSq2dA4gwUrK04Xk0+JpkRP1kG40Mqh
vYTvUgl3yYeHRgjT+Okl/X0T7xeyD/S3oxGSJ+7vJUBgA6D5FiJ6+RTLM31WsHnm2/dGpQLMYqgz
vcXbI0G+kHwIWh8r1bHhqcgLBlNJfFNvRG+pwkkEGYUd/MBv3/3oS1JOd5gYxRkPa2B3pNyOx07Z
T9l2rNqN8GQqhLghEfK+D0cbTEwsnft34sHgqPdeNC0UUpSAqEb9AzihQ2ht9L0OVcb/nB/xyMkF
unuU/7Rq7PPU6NC/6dWP7AV+/3u46J/POxtdFKCAs1djmDMfQwC2NTI42dQoxqBoU8wGjSXXg1k5
Bl16TcdVFh2me2dfJhuQI6XKT7wJ0Xwh4rwIlKDFy9gE6iK2cpa5v0bOoFn4c2xdCAoNoKY8x3mJ
mcYQG5kpi4TMwhvHKe+TtCJOA0Ss9B0joXIrKkTiTNPiOTsHkQpjuXxSm0rKtD7njf1OdIY02wyO
M94gssIwqW42o7D/nq60arOdz5MoG6DgUIWJL1VH/60cO4crzcNcH8bpfLakNTJSOwoaH0dm7X+o
IMRWMMOywsDxa3r58gJYwVorzEANCwvr9Y7xjBd4ZApAwQ5Kn/Xv+3t9TKR8zXPkAcOcJxB0/p5e
GoDXl0gH0UGSlPpO7z1dy+fWdcvZXSa9XBv7vn4S3CK07+lxH8nbcOmbgwV4jYgcrvULC0MjAlyS
xOFOseKpsXmF4Hjq7Z1zjiL4Dceac73rHdINV3cie/k36pOWwP5VX+QxiSNWJTnCKrXaXxqqlM0T
T1P8CSwivmOvUHwkRF8hlYu7ZGYvbZMf1kimWuEwctsudbU5iUF/hsIp4PaiF0IWjglVvcPS7IOR
6zXdDwPhr49vzRKw6/hp4l93A7yBBFuEl089nC3g2rV9F8S90y4PY5YTUP/f9GmVqGnESegSTTHW
lKznEYJToLQNak1fduHWIlSb8+TjJ/QQYdWQCTpv4rAXUZ/iA5LGKsskcKF8mPYnW+fl1BLRscmv
eWHuHEpxwUozDTVnAjlic/WfX2fGHcJr/7xFIn69rJ37LvPyn3ayHmqyTKMoKPZYnFrjqLgSQ7X0
9CrccvzLuchPULbBSYjkSoG3hufobpwGZCi/SJ48eETxh8nQpEOq7AsCbdw+GHx1XqcpEpk7ACa9
1IuEke5ljQ5zNn0qpnyKfcfXZuGK39NS/sP7+vKrgO1tkAy7Kh9GlaDPRQQcORrpqlyOhP6f8nQG
yO/7tOGijnAeO1H1ZbH4K8UIZNwPBRLAfHWPNfE6opWtfkoIrwK+0jlYz6WMCjt99qojFGEhqoGf
2NS2xbroofJ6kvo6BOlT+EbG7moSYA+0jxPrJydnOjv6mrkCLR03O1SsP+3mSZqMIvR/SBSDPgjP
X9PPVlHIItSIq87ELKMVQuGyg4LtiB1U1xakBNWpMbIAo1N/rE5kSEw0Bltru9VeayE7XG6+IQZI
PVh41WuzncRQ4IoTOR8jJtrjA8ibV4xGvDpTgUK8UaG/DHn9dthXAZq5Qv4Hpb7QTbir4W3HwPCL
qZja2jnUTUmxFlDOiF17xk6ysP/MKE5DvyCVTIxZrOQuE9YIGegB8U3fraVNEP2uRY9npLXIb+a0
6DnqDg9ys2UVNmMg3d4iRB2AYGFV66XRGNnTjOZap+nsxj/3wwMeExIVmh5IH8JN64YrdDDjox5e
0c1UE8ZD2p4e+Tqd2wqW0tMNKnRj3S8jDODVTU5nrCNMAJTKHQlw1xDQRRkpSaltIAA2NkR+MRFG
oWVZlc/TIWENbPkVfc5cfQxHfbS0bqps8HS+K8QgpqUoSD6jo9+Hcv96SLDNGqV/Is/w9YmeZYA8
CI66sS1Tq9rvPTYmXZtpshsQJEPzBNguRSSCSt15yShVd236Hgvu3+oioz2CN1QHYNydBZ03OQ4D
qXl6Btv47hOUZekIrDlhHuQNgL9R2kRvFmOYRFtrjyZGFnQ6Swza19SQn8sRHw66JFbsnefNblc7
FnBJpGcF2fQ1s3rnkgMnA2Lf0FkkqVfF/BXo+cbd15TJkTCxR5k5GqWna0qk+nA1eyr0DlRSzb5d
ayzLaema/IDQPlQ8ZZ0S6LOfg9KIg9EUj4i3GdTuo++uY8aizm0a2vPLitn/2ggI7r/5xP0CgEbB
Bu6Y2i0tAbvdubHmiFXMFz0hqkHBMToFvhv4YjoS9Vi7tKUPD7vMZ27TwTe6IiP5JuWr/qZV2V6G
85Cr6jZGOc+VqJsXuj8gdQfgqCJoyNxk8xfcDZL1kn9rfbFqE+tQQr98vuld2ujiq4JrVVxMS8OT
AFsvddNGOg20eaaUiABYSRss4oFxtmzBd4r4HKbpF8RyljsgRCp68vDSIopW0oB5Zp5++I0iJiUM
P6pNBRRwj4RncfIDWNLhv3UgOeXwE0UwvFicvTKiR3P+k4277tD0c4Mtionr8HwPst70TPI/bSqz
mPDWXKpmxSlTnilp/w3NnB3q6EVYIbCwA0nxuXiup8zByN3cWy1wf8I2w9VnP7fPoeSpiuOrvPuy
1MVE7hcS5q/425yWK2f2k9SOHaXnRdrB5jaURFy7nLV6S1LnyHFH0i2zKU0TkEutdC+7TIVufynj
jdtZlRlCj33MLUfs2j5Ep5rjLp/jBv9HBvvyg24uMX5pinmyYfOKJUvvBzoz45mOeglojWWVW0ml
FRjLxonq5LDjm/RYWt7cFWVrepv8Lbp4FbokTNoVYlE5x1HTWVd8pOL7gO4brOHeiFk6jr5VT3b5
h/3n7ECuDvmPxNpMJto/a0cCWPPU8SW5Kep4n+Z2a9dGGBJJdG9qUk1FRi70USn2ii1NllcXhBIC
s4SLOiY7EoQtA6vD0vgCOs5Fbo3hq+K+8VaGX8cyOfToxl1EEhcDdEAwAGynfFwqGMNdn0euR2/m
zrPqClu5RGV5rZ76a0+k3+HeuGqE9sFAUrj971L96PySxSJ0QegM2KMAbwM6x+7HXvAN8r9B1t78
GeCks+NNLChyNKQESiLMY+zJIhlA6xp8Ye0190xkHKWC2qTRJMyLQVfXEKXMhOPDDclqLM9wt4z4
kiVuhY4XeZLhV7EvkWtMA744n2bAmjuFu/+ctIy3bOduAfCKCJCGjT703I34/wF7oWpOJzBWApHT
gyBOIUhDPm1y2rg3y6WhvZfQzPtZldsf+xnQs5FUGhPnWEGBUL7XZJOEIbEO+XmRF4rWQfQC4t7C
x1HJPwbQAjsEkOyxAlWvtiT8/OTqqIuy5EtmYwW/O1uoizMvi4SJdzTtU6YTkHJ6dFrQnrWoarVY
Bv84i2KTGg7k5MdRrz5syOeIwZ7GnVm4zoOIDHY2/O+jffsU7UhDJEhLzgDAGbtYCktErvVTszOQ
7Ms92eehpZiKC3JVMfUmvtIz7cscIldrdjxvSEcV7AokDsFfz8m2Ln/kf0xJUSiooOONq8oZGkd+
cUXA7i7R1BJS/XBsruFUK/MJoitX51PbP3OuYy2ZV8PADBfoICevXXomOTd3+BrfYOXaIWRbAG6z
glNO2gTcEcD9wHkZeVCZy2rI3gbjhPfH4YkFIwAm2OAL77EfCmyhueelezAGAqdQ29aTPibthxDp
l4soq5pL2sTLhA3LNAyMiIIZBV88wWKHxU73iigQMd9G2+SA55X1X/pQXzInbILajuYVEQ0tHpi7
z49u59ooODnB6Dk4hyJTZEUqoJu5QYoxf97Ob9DJ2DrP5fQlOT+J4cIYqGY14Cg9gJ3j3K7PU5Io
zOpuoRvx/nBMIM1eeWUSzXGFkfl61movndKB2AlhSFky93ddM3PRP2FgBr12fCbPU8bpr2innan6
kSi4BRLP1zhKeFmEHT0PYmouzLJ864SQlrTvS1whpezs0zoS17pNKS4zrxZwwqc8L+9UNL9P1WGg
eL9g+b1BnzMbGPK33Tk/hJ+vIKx/OqGQZfp+sA2GPYncM8kfnBTIitP6RAueRF+iN+W0j//WyCpI
O9anPbXnhH0fsf11rdDpAGkAUQOpBJd2GnZs5GpocV1kEHXC0i8YLg4SdD2PBheeNxr9q7sv2HHr
INZD3mkXeg8HLFaxhDazkipFfhF97bzAbdyItOHAztcF74wQo4z+pqn+9uWWOpNm3FKX+NRazRX8
Eg3vlgh+3UhHYwejJ1BwwfhMVvX5Wh0wpBODziJxdVSLTAvnnCe+KagU3yujuyoma9zF3IPowYB6
Cj246yAhiJ5Pyf0TDXlgx0nMZDmCNiq0KrVrGXSZPgj2se/2XSHm3MVURIg3TQkHdFvHuUTts9ve
oL4LUrsbWiMtLAAQVrtE+mKI6hvOFuALr5QeeCRogtX0e0uESIuf0jzjWOBgb6d3rTu1zH2S6Nzn
VbAcYD8pvrTE61xilxt/g/xGu85JTXqMnTYpJB9RhRoqU0V6kV5vvoV5VzRF5PgcT+7KIqyklVx0
jZmao+Xw3ubQDbBQ3birFhUr3lLT2BUb5kfc1h6H54ypAP+8rkmjdJ/vicfCUDJRgSManayu6/B2
j8hfkF/kC+E+XIRZp+Wd/Bv3usWjec++uE3cXUaZfnQ4SwpnP0Xj/L1b7Rt1xWs0iihLcrZcn6sZ
LsaK63EILaGwZx0mOQOIYM2WhZdHUSt4Ka2qqvDbXTy/yodiYu4P6iwSaQk68sxMAAvl7Hnri4K/
1b1WyU0KNOcvEhiTiNZuXbe74qaWW7lHIE5L3RngB/Upm3Rs66JCDcUgS/4Nadzc0z276U2WwsKw
5bA5mP9pe3+FwjkQH5JuvJUd60ogPBDBVsyD3rN/5ZRxm56Dyv5Ax8T8UloLkA2q/1cUfXb3MbCS
HKW7MIs2VJdbmfoEr/TWe9MJT66XDEAlvMLbP8wR8KWz5tbg/lAMSU1uX662KxasTUPUq3uawrEG
GPxRRzUcHOTiAQg9aWBvq3nZreJ9crENlcKIVUI2VgyKicyD3vAQvHQEIxRny6e/cc1AUnWs2cpq
swvI2VfO8bj56ATLMP4QlHf+E9VUc0bhyh0gI7cugyzDFBJZ5bYKisP878THKk21TlCPMrYaaFja
57hA+RodMw+WMb65SQdCztdRiemMlYm8s/xjz4WM/39ah4GU6cwfhHFvVBfiNdr7l3v5nqmB9NZh
8akCEMP9K4O16GrBXTeNjuJ5QG2Pq1/+a64q256c58i6k4SAmMfWzPgUrNbyj8AJZVtRR2RseBzM
d7dioUFo37d538thXnSL4HUTaHIggrZZFQQ/NtK6qfoJSMCGc/zSKag8Gu8qayY0dFzHSQuAlOZC
/S5wdaI2AmcsSbnOqMEmKjuEDVaznbZCYa7ZXUG2jYbJ6d4LmlRzqjPbd4MAg9NgOpKLtfEFWCOt
LkFReOjYZSDGnH7t0uxDUOVMPgF7fg2ZzaOA2xe32CVjB7tIJnZjVwWM+t510ttblcqn7BVqjnq0
G68akMTRmCnP3sl5WTTAlcFIWna+dejYLus/fK/XdlIeDbhaMpzNvVy/+eLtWyIdiwRF7LOXXGq/
Z9QFgUlG8fShMHIqjkw07po/T3ssFKeqUgObaYOHr8IUGSZdsFn3sPfatm4awotLl3omv1c/z4AB
EZ8TLrWx6/lA68GVY/TQwMYSbtQTATqULzambk+h4cC0dTJDY3L1KGrgONAJdx/bP1si0K8M1NDk
FjkfUeJ+eyZGdjPDMOquMWLaNlk3jfQ2kWgxPDVkjZlQIu0aFxQnwyLlYjzxSr3zpINCVdKhq7L/
4NdwOVG3MYlCsc/RJ6xN/qiqhhloRNL0TgGPmwr7giXHR9LU9/pnn80tCGJBQyExw4WZoNMLDygG
SOeQ7Ai6fa+JYBl6YSjZgBWxRcaEZMxO0fPkOkjJ6uDEhORiCLBIk842O68/qK07/43LdY90OUld
oYTQ/beOJ9RR7XF8EPcA850Zo3r2cyTGZC4ilN1ep6vRKdEAR/3Q4Rf/zEvMOQ9/83NjBA8cJHfr
t8Swe018rZnPk/Fa7BYA1nGsSFCON3Mqmy4o3dSt+nc/99N4HlgT+iRoy5yt12FixueRVP+ZLJfU
L3Nd7u3PIN3RgC3M3Fkt4OYLSAyW6bsUgxO0XBmJ+NnXCI8HH/i3z7kJ03YUsE+92tpZwDhVc1Gl
fH9efM2R/BpatO7mPOz/QCSz7L6xIpBSfOln6ccjewrDNhfY8GwGE1wLRp+8HuSgtxNN00LT1AWB
2UQlpRSP6o0cBkgu9zbLCAie8zEaj+O6g+C3L08cKiZ1XDq9Gv0NpYVjP1tD3WvPLnFeSfOAiCez
6eNPl0LX14qt160mm0wbZ7c4c21aZQM/s7k569rhdw030p17rjQ3z0cW6nPImAhmpoPXt/1Byyzs
kiCxVzBddqFwVbFJqDOEEWB65DiWibqpSykzWdfbZMpktOFxsS7RY0zuX6jIGy3s9kYulG2sjkOE
+Zz6MP3WEBcs9Uq3kpxQxkVb2M3LKwab5ncJYxLTQ/JrjIr8hE99sPscs0MlqCQubs0Lft8iMmSW
EaJPuIcv4cVT5Ty54Ntt99XdG/Z1ZS9eeaog36iO3enTy75FhS3TGylWIf54xrgSx22MrjkP1Kto
AhRL1ZxFM6bJKk2aBGRcsLA6mPQXl24U5fwPiHJWGCH1zRmnbUIj73tYJbNohaC0iwu7xYVR93WC
SeTpiTA8BpeEtmiNi3cZPsxtzSIC71wRS2DOssDodoh0dJNY2DOR9+4/FCV1AnKr+sumgai/mWyd
4omBAHVxxbSp6GaOwdWh/GYOCazA2oocwYLCE++EdKIxwL+YuecVyHDDtapuHaCSt1GcSEvIYOw3
AjZmUwrpQtNqQ4npi8rOVbuCzYIit1uQS/msmRXteNdFIEPNpopYlPYDhj5BaHtBbiysDE0cIqTi
ZzZJR6L00FV/TvKOWzws0VM89sId7MpP4kKG91pHPyQaIOUlfEmZTl15Fgk74raIgCkscr7ThWET
WcISrMz/ivr/n0JEM/KIVo3dwO5OOAiYagHnJTjhNyePWZy+aOLq0dLDCl+ErSvhsfKVsee0eujT
CI/5r/3qjxo5efY+MwktKgfgdfYdgrpF23ifFf4uhA7rea4x4emyksCePzKQJNzDcxtu1iH+uvNT
kxSueUeJ1Y5pbF1CIrOmuyjCWzU+AVaea4nsW8YxnONNPkMuEVpOBUqscLCgKwRwFN5b3IdaH86i
2NeR0Wc8l/lDaeVGBZROVo0QLZ3eOMLseq1SfECvUVWwyDMpJeUGKNAo7V7hujyRz441q19noRdM
H3jXdgLnu7DSOjS0H/eZ2XL+o6rYbF6ZtTm37RSSY/Q+Kkpik2YwHOrf2fECmhjdP9R4G5pdCWOJ
WiTWr/Lay1X5v1mUJLPdrAcY8nNKO+xb074uQLXIl5uOgfzYKqk90ow908MneABhOFa0mn9O/K8k
xuhW0XL5YOjQbZbXuVkbRCOz1FrC/PeFWzQTqQMSqd1c/o7SzYW3f3VCjo1Yh0MYh4tZeGDrunw9
Sy3L3UZEkqn+ZdLqB4hWqXtIN5r/GP+qoHHP91YmJ01bvfdYI4myP5rDsqZy+/duSu6vfVh9NSsC
Ejx8W25Kgiz0B16s0wbpB/BLLalYjl/eppy3Yhi56soLdRYqp6ziJz7dOHje/3V8b6bABz+97Koh
wXfW96t7cDo1uGkk6hAlqhcj6lIw9HhpwnGrjdbcRDVE3PWRtdxNJF3NqmDShgN4OWYG61RcwhFr
QFd91ztmJpccm1FW0UwaOvQie61T4ujhn0++dyYJuj1/WbK92rEt89AIMquByy1aBvloE41sLzGT
UiSKTSIWFHFk+k2DovKF0jKSBYTd3y4gH279JLCL0I0XLvs1bFYDivv/isgfux5xPJavLnpbi4+I
DeS3Xuikk/9iqCDSImilkIBzw9S4NftsGbUpqy4sY4L4n322njt5czworWI2rG5ExcTZoOORHEpo
I9oYkISgNss/yF11+sLwa3+85hOmPdnPITq0Dv8QfkXUeMprRswzbBdsPrv/+NH/kzZnGMkbf3Hl
/9RxPuNnK28q1Mm92wOYEXKGQExVe9yua/mn8KU6aEgZFXLOoA77iL+1p9+fzMw01CwqeHQspYr6
6u3cmOxyqKlEJYxIFD+sUWEC6q/w9TNQAYS2GE1Ft3QMi87uMr6X5d3N8ABnj++Aim6msO7R2EkG
JSFmLyDUTDvSWLWJFbxmKpT9zIt3gEUnL4hTsURD1n+DzZM8fr0KN5uHWQEe/UPKIecZaYj0oe96
JG+0XSPH/BdH0VPi0xboS7Kh5ts8VYCNh8DtHmARonPl2qtXYFENLwzLOEdWN1nlL9nNOvhVfAxL
+zBUYl1da66vnnT4u9rbPMspt83NjSXImc6f82awZuYjvZ1oO98ZIUXXFHsq++2z7mq39gtTCpul
Q49ZvvmRKQqd3Wpk44E9c+Lv9gJR4EJCUffi/FDB1gdQoRqfib1i5cmVapBh2E7P1L+iWkeeOQeM
8qS8kQxg+8XjTMoNDmjmwe2qk75MPDebZaXGD4q462m4NTDiUBmtLPVcBhuTcMMqyE+MB3Lr9FGZ
PCxZ5cYeREfvLxA7AGdyAIqX5356eZ0WrfPGpAedWef6GMKHZPzupZ6EBy1lVopRkWWBTfyrNmws
Mojl6CgHMdWsu6jqPK/boBGOEbHPoEnvN58SJegGDKxgTYg8UVcgCy/utjIQiSL4dJ0H4LMTkwlb
foCYQtQ5MnFO/R4FHoftmaXjR2Ig9v2WzqP5p3M8az59tExEer/WXJyd4Xrj6V2KzWoSrT5K2eW3
Rg5lESU9BOiSTiKi9/DpUIEy/VDqQIs0CGQnH52DZRyx/nclz1m9t9b0SlfS17eh5QY343Fw9q4c
XCl5kofQUjlao80Z6gAmBxjMRarpTvLzx2XifL4HRg++3+dAxIyqD392SLkoXoU7r+fbCye/S7Ya
5nLHQCucNluAidw9Fe5F7hOJGbwJyjbr0NGQ5l2XdHSkY1PcdX/w4icBSVWkeF8F1JMy5MFsYVyV
N1R1JSBaCepTk04O4sxqwrpmav98pfT06xsFraHtJ/6tDFfHuOxYIgGOO845lsyjXCU6tglVVWMy
LkJ8EOYfYGPUbokK2iH2UaK0r+DPava2hHw79LrE/kE1Jpe4yWST5Zu+63EOpMOfoKf77CdYmGfA
5OmrgHto8rHdCf6atUUSd2E85GHKJr+hvXoo7LLDhD6FG02yjS4wZaoYmJtk/mjGW6G81CyWHxM7
A9Rs3+06cMXp6HNdmpcge2CaKqNM+EQoqJZh6uNjNEkBTgJV+fLP7m+XNdvXQvVsVqX9WIlGSHGi
H5skELHDPIjIR4Z5Bd1euBvXbjoBDIgeW02BzbmsGWuW7lkl6OOdOYkfabV3fYvDt3u1gD32+qA3
pUcZAxPrmOOBi8HVjpXyhwyJHy1YreK80kv/ZXEXFZRqXEJ/JyoWhMZiYci7bTnCaCJM+hpUN6Nj
0saK8ywv9ycYRKZ8JK1QLmr290gIef8A9E5dfzUkRGwT/An+zZYheMXBr26eZbks9mHeQy3pGC8e
ZfKUt1UASq1JbmUFYD0Uae8px5gY4bGmTAvcrfMc5oEI0nv5dX/cIAloqhwkhF0s31/aDXi7C6yc
RVmJlpNAFiCCUbgTR20eodDNPzBBB/Qk+gZW2i0P5I7A052q/quUtTmNEhOYSV8WmYIM2m9NzWQ0
KaB8qh9cCbC11wRNvfW0Vw1youjknwId+M7WToz7K6A2Kgy4qJ3ucpKhyQvwx/OSHZVnkpEYLgf6
1BnjdJQTr08HJC3uvD5ecjP7ajSQtS0K8gnA7ql4k4zkSjWp4ONiM058gplEowUf2KQ/ABZdF2Vq
I2NKsobMS3EvRy/8ppQ8o0kYS/BqiSZ1/mJz5ONuOp3tihBmAoZjc7yqcH9jDRR/CmPO/Kbykzsi
WILviRSeNXHvj17qhEDGyJ/MpdBLatkxAF8q9ZfM59wSS2mkzJVgKmxDmlYOk9WgMMxfiyp56bQ6
xJQ0Cn1aHRUitvirpXhQUmLbHNzchQpVVfYinrSD+9+V0jYslVk10GWcNqx/G18LQ+hQAIiLgqYc
FUQk/FXgSxJyu2inzWQ01LtxBx4FnK6fkJKr3eQv6/nbF44vJNWECGsTmrOv8/Bj0ij4kEQE6yk7
OWIqEMnJvz48wvnE9stTtVoyd9zRQw02pChdVpqrjqF0vVG8U7uVS35Dt4XQW3SxB0F3GgRjIXfP
Ccld7tTX3MjE1Lfo4kfGfEKNgzzQdQMI5mAN3yXXaog65dF2YK3C/Xo/XaOZLB/JTiA2cTdwHuzT
/pLyKd33U3u2vIQM6l1djAfZ8p0QPAyHWehPp/rat+0tZuJB+A6WbaNbeSuPXptbiJ1JeYG1IgEk
yA3MlCQYvE0OmI8h3tBx9qo/K0V7um1ZMtgOaG2ZMCwpWiUiyLm8MfjNMUXRz1CoF6FLlu6gsSmk
WPqvohm5FVBjjm1HM9nIYr17VAiK05Qs+sxvPqXakXt36veHST6lWhK9eB/2JuuN1Ueg/aDGv7MG
1pwpZJLOLNxokEgo2tKCRyv6tS9pQ5geYm/5RPOnw25s4gawyLU6OnnM1vPCVORXBwWmvy9HPm37
csMn1R39M6XMNchHHU5il3Fm3rD+evgdeS9M1wl54pIBbEdC9lthRIUvZkrPvb/BZf3Qbncbq0n4
TsshlEZ5YQCMTw68CTr3IUu+dDTmGMlYgenbH/422XT6xXkXveHJVXrLX3uM1RfMH4E06/NC22aJ
1GUiDG5hNUdZTN6bY+oYBKCrrEJQTA929bI3T2YH23x1TSp3bq3P3OtZBjrSP46EbZDWJgwNb6f3
pIU0yjoxjuLS+ctg86+UAME45BmFwp8c7rG49ZBzs4d+zBrjVZpTJoZUaVNT6O4BlWQMBdYNWRt5
SuxVcRzM6liJYwYh0IMc1EX7BLQXStLzsy2C8v7ZDxtonhszIs/LF3z3uCNvnsYUHlw4h7mdqj+s
WbRkLLvnae/fE+OJMP5iAPBf+YxcQgANWKznGIS8crYIKfvERd2PXqRwe7ltsySXksyPrhlF7pvP
YicGeKMcJHY2ExfMcKl/fnsD7ULqpf8wmgBuxwJWlheNgPMRLFLBM1A1VemMDalLoAcsho5AQ9Zw
9vjU2z1g8JfxQXF/cyXfCdm1ncNWcIUHhbMbUoLxP9/rC6r+XXKt1tNEFVmGgDp1sG9HN6pPPNrD
bwZe8mN8jqRCd/IAGgFeEH17Y5Q13PPu4+6MGAGW3x4/3KE3c5Rt///OSzZye3/Dnavpm+GqRXQP
b3evLIm7qrbTIREfJ1P7tDmQ7qXiAplk6proQiZasrhtAh4WbTZuLXJT6DMsD1aw67e65BveDUkp
YzrHSsNTDB0aUNi7xk2emtqyJgj3sMatLoRuSSJ4/AO2bdTFLh5l7mXRvRN6NrXlLq2ETYMN8OQm
yIVUrU26xia8wqFY2yWI3ytpeM7yqRvmLOtxwVOCR5VzJ8/ihq7SOz6PfdLSPOOu5xtRlWTXQRI0
Typ+a6u3SXwmCnkbRQuQWqGNG/WytAUgJggCh5I7TK3CRPq+uPVU7m9Gxh+CmbxP8iGmi9+bxzuN
cPcEDyVH9HNLPGGfquGWuM78xMBjGAUu6WrCXEFVLTjefv8BeySZPZ0o8egHCjBfIOyGIlH+KSbH
mVsqz5hfuXXNBnXgcaeRPWp1toRch8JXRdILiBxgnJLRMPAaXxjws2nmQGWFJ9e7YAiTKaQ+O5BK
Hkm9zM73GG2SCTLGb/s1qmqZeqhJDE9yCq/jTr9RexW5snJtE61s94MAyDZqpepd6tYE60DVaEmj
+eORafAyC1mUxymYvDx7WzHz4yRo1AsnFJYTFL+C3e+g3Fa9JDyoDBUm5LzfvDB8R5/eJcNeUfnx
KxQfp40bR6Nf4kXKVAYWMRaShMjHhC5gmfnnXhOI5rkGVD2aM3c2ipq5gQiPi2d6uaFrZ28QANk9
AdynkHddAhzhXemdyDO3qGPP0V0bSrsN5kapUuKkOjeOZv6DBZ/YM0HMJnusYrA0Gy/zSy/WfmTP
HRxEozZjLko+bA9ze0f00I0XC78u5LBvRaCXa5/ADNydhk4VWUHX/g+G7XPQ0joYhD8pQm78snJp
TQtsYn7EPfvMjqLpogNIX9moZdcQGHYQ7wGXsQoJwLpa6Ex5/zisnPU4GfrR6AAO/HLCQBJ5uKEK
vSqrWmMOhgqns4XI3237j3jcr9DRuQjeb5x5XUVvsWatOb8VI8ihFxxK9PBFOJ/9HlecsxtyGoeV
9FS0g4fvHotc/rkbN6fNP1mLZ7fzHmc9Begr4nIIFtOg6HObikPL05gfbaHh9OTM1CJcotQGLMtC
7B9f6/6nORXdK+G2vWRBukPKERwdpDWkRNUkY+esfQ6YVyFvTqJZApANffGf5xem08kuh9mxFgsn
E+y8nnTWbkr/3Dvube8pGqUGfWow9oTQcV1PP6N+HGriigvxr4iEceNZJE4zuGgie69vtK5igLBo
KsP/izBqAIx5R8eguXDWYNNPYl0KmGNSWNSs+8fm8GvuITjiUJpC6EZRF6oaLdaieSqC8DMNdAkF
dfwvg1TtUdujfQIqegyRn8027CTxlpdN751M9vkui/jj9cZNnY1NxYZadvZMGVYplOpRlkLYHGHy
NyXuDZGtm0YviVa6HVsLVfJnn01g8/gJPBtH6WeVmsVk2DsqZE3it0yjuIgkLa0XM+053WyilsNa
Y9aCG1h01u8EoLNvgxoJqj1vPJG2d8sSTfCezfrQITaTzlji9/IsGr0DMYAGaoOTWfSEgK1mdQWI
rlNYvS+/zc2zHOq6HjIvtkiYJjNmW7T/gyxSe/dGTUznYCOR8FIjXWNUv3v/GKgS6D1fbBIpqivB
zLHr656o8J5BCQPUFt7MkpR4RcvYoMu/9UWycJn+/37vzssq7cqhEJVxptBgyP9Jv/u+L5Ubu5vw
6dJJ5UoqHmLT8w4P7bhrOWxKFVM3RHK+W8THWz1h/ugWOVoy48B5Ch3G0KDmofa8Sx4pul3ES0Zk
bxN+fXOBs+/YyfEV87sU2gJ+DNEdyAQ9C4FVe/5nQ7LkF1SwGuRXXmyeT9aIELT9klLtEDn48hhm
gZ6TN6G/apTHYipTKAPlGq+10+kH7YAs2kSLANOp6W5rXCP3k5yhTYXce+ohnNZjr/GIQDjdq/0c
jWUptRrO79WQUJ382dDzfwSVwUIs8lPv/6JTCAoliJRAAO9sEEomEseGb5pBR710G8aAl1x0Wjz8
WfG++iclTEXO/2e3AcrEoPdMIMIbnU+L2Ez8GDHcLMOEApwknKhacl17UiVDHMcRTzSJ2Hz46PJX
iDHnfkZ8bivyerG3U4Ywa56CDqjhNbdQg35siCnhMQJIhRvgBANLtPomdNHXEIVi36WG2ztPtk9R
q3cKnQp+QzCilwFZS+A3gxlwE8ZGf6JI1en/XmIDCvzmx80uVVOk/PeFrGB3sPV8CELXfGA7tpJ5
6Y00aKxfdpAwpe98J0bT6d06jH1W3dvN8VWFG+wITlneVaQQNF+zB0xOTbp5rgoj513n/L7Y8rbk
chs5Z6ZF6hnkympXHVgywIHvveQw7rgH2NSx+V/D7Qo3fiToS7UMFQQjMJ32Le/TTyHQRvn9Xg3R
JtPK6vAYeo8rObwMckvxCjaLxsNbRzCCjzA9tbvisLH+2oIC6/dPq5xT3fSICGul79yI20889SOP
pUdW9rMu66WXmb9+bIkE4eh4FRH0cXU9rYv3p9YnuDMBAlEbEM4p2k2HFjL6Mgc8MoQUHkWz4zX2
Ahyh1FeMjfIyGwydDUOqFXMAEBUrnHznhjPmKQPIQI1rgzPV/u1cXS9GsxdWRHtjF3sXjn5Du96A
IdsXhMpnKgozf6VS3gDrFrWYOfyEUrJHa3axBv+5CkUaP6Ovnt7D7O/oOnIso3QyZwsh/inuPxxf
m6PUNdOPUEiD2vbHEUZwzA6jcvXhpFXQkDd3Ulx2pul2gj+Zi3JHiv31DFRX2YbQJ5SPqTIKIXqW
n7Uhx0N1l1bQTCGuc1646AY4F4QgpEe4+0UmZHW3oqCNN3ejEbbLxtBrMmn3vtlfGwVeGHnqlbth
wLmCmWekX+1EYeAQiqx7+2oxsaRvi0Uubsto6TWvJyWXcq81NScHGc+AKFaSK7tUlFrWfJ5alguu
UxiQpUuPz92zBkFrCeVpLxEI4rhesU4rP7SPYkJkoy5nh8nBzr+4Tz88JyKuvdCWMjfczZIq8a6U
Km9hhV3PvXyHCVzQm5h4F15kGxu4KI6ldq9je/VoebnVh4As04OlP4xwfYxb7svKc+YkKSEy2IA/
EElrX0h5wFgfZ7RddcxwbMKtAqNVLRQOQGCokW1TPL8ncTwCMojHm7Boqgs+WlRK3wYaN7iCuetM
tjOdityT9KRBZxKnLk2Be+JV3NqkRaOLwLXOPLTbPm0N4aLxGNxWdfV1272xJ02KWZBxTCuMC6Nc
dBymCy3WrS3RSEQveq/dWqi5s/IJmr5lxTL0u5t3qgwtIlGLEv24YC9Arw8EIECbnshmwbI7hIjS
Y3XMth4bsFFroST3w80ig2vph0rWRCn3yIGVHi+bmhGR6I3xwYfSmyjM6ss3c04imfRmUdu+L+aD
EU1rFXyxvPzoqdi2LYx75tg32kFZ6Y/qsd3AvgD2oLaaN27t0zJotM3vcsTxx4TnThSsEZrkDV7A
HfLk4n5cHrc6vJcgQWZvBevEopKYHLlMHVTIc3pGilGz8idIvV+sFCUDZFOlYBAsyZDB1x+KlKXw
71JAvyLCwUts5ts0Z1WjSKL+6N79xePHIl6TLtSOQ5c0VRYeksXa1fHD/5phdkqA36ih6QuAHESZ
HHpf9IgaHXXj0CUyOhvJd7iVziGd7pjjh/WEq0V/a2/Dwb7sdGGJ2iijr04rZ78Wlb/oY82E7YAR
NVI/2gCnvviARm6e3tDEcRgtqeKR1WCaLV7DoUCFJlgCz7zZTZVC3cbgfm9c0r2kZmiF+yska+kt
5wK/eidpIQsVdHwJjyATe8lY0d8Cz8jkcatUIGcynZdj08FSpgQ1ovQRsR7tq7sVxNTzsmSdU8ZC
DrvlMLhNKFNwmkdGYko7TJjFt6DniAgB0+v2xnT+OYidFpfZz5IHirjpner1VM/+s27RJSH612wU
tjJ033IhMG7pjdgMr2AiTjE3r5LqQIFX/tP41Z5uWP/Ug+wXt2YCPdSsQfQK2hABo2ghpRdUVDzB
hBSYmU3Sm1eUJeIvz0kTlbI0syC8BgU6nNPuX6g4ZqjGP7FqEzgvgPleFm1RgTBa7mLmPLgplpZf
N08TO52LO7lCVAtUuJe5hB5JyKDWlCg6Xh83AybdUfKCQFp8G+6KxgGD0RHjHFxcqJFW32Na3LOe
yBc+rNzMXH8YoO6q5gAw/3gTtXouH1SXt7UlCYV/fep+uaoHmvhtMak3/w0zn9zansTnOdFIF9X2
2ZipKBsB4jjE3qcVhUcFusLBpPkhIYqK3UP2Sw8Xy+0uiJN5Tr0Nnyc3Fqwh3etkHUV1UhRRiRME
Tns9A+Nu4DcPtxUdq1jeKaHtUrAyC+7QUQWlI87ZV9RuyCuJStd11zOeNe/jBQ4aftlEP83hl607
uXcLMI+sj+98kfYGfy9EtBjpX1FvMIkoc2TkDaVSgoeYfDo932ghZU1tXumxOWglzTYua08lFity
yhTE9RQdkEKMfpFh5A8PuKeNLZWxkxHlxRUMRUTgr5Jrzzj9V450ReXt5+nfi/FEIj22TQupF65h
MRDfTd/tKIELwxwq/QSVzniUS2AX9bcIV0H/i+jGKvwu4NvcJXnvm6ie4MjppF7v/CAsxii7UvrM
NLu+TnLf26/BP2SBDIAWjrg6fm0lusRVFC+k6EsptCEoC85/Jx2CqBnfpBccBzs2lNWGAI3x25d4
bUXUCnoFP6XGn+ZXBT25TdQ0WvL8pU2P+M56R+DwWPZcGJMZWDndt9bFepH5JEOrepk/B/ThL4QS
Z4s8PcKtU9ouDEdms6WKAuZEn4K0QtgKUHHw+OWkm8HC5rcqO6tmJ8iKnjCIhDbpZjI88ODyV8vs
c9UZ2lSnh0TuOsTr5HUXUOErnnKL2IAf0I10VilkvTceSgQ85WWuPG1psUT4VcGYABRGm7ZkxzaP
HIoqRo2pPp1LLrWE67iCTLX8/OftEWC67bUsdtjPYUgSfZuRNXKfdOPGW9/bROlkrjAyQKff5vXP
DJytHtXoi5kDepAZNiwy8A8Qzdu7tIcWo6NTAIi0sVV/pd9L/vnkxvFqEA5657YnIVLW+QpAcI6O
SEMlNfZ9dAehRnMU5ORrVnqYLazW5JRfpq0IcOy/eJK8mEmLXL4fN2RCW8FOOC+uO3AAt26yubJR
ZmpheeDF1DlISeEZJ67gTXzHEhbmqPqhhiMUcRRtVgEHh7e6kAZo9r92+Y8QCiu804apUlayqQJG
oYHd8DdcIe79aXBNH9+JnXRSORckW8mf0GkRNJb8TfgODAf7aNCcVqjA7PoKXXLt0tzzis+Cd1bG
XmTwEQQjGwGplyGovLdhE6ap8kI9xQphzU8dRUOjtJpw3rxL6m8UDmlLdX/e+YujOkYDK3Z2eGsZ
wX7bSFxQnu1TLVBOo1KUExQ/fYzNfAdzlB+/+MVR6k8es8yv3p6gZGSwPhHgl+GqtFeExz/kColT
YgJrjEF6Bt8WewZshAJMpS/UFaw9GaVRvjoYZr2OXm7jobYTCYwcMJ1j1Dcy5ReuSkEelvSPDhpf
Tvwr+sNd9RHxHULXGV6fLNbeUHdEuBDhHbnWzO9IiJqNXI88n8c3vgyJw8H+E6fSCDD4Klh6TjI7
LoBQ/WBIfAOloIt8oFmCXiILVHDRqiP6q1Q9JleoZa2lDdEME1thkCyyr9ByxZog4LvSPv8Qv+CJ
3qeHAcazYtLw5wwBgD847k5h6E4Ow7e6AjSS3PPpE0GRcmi7f1mEx1bchMrKxN2oijRDgiMbgKiR
BrZkQ9nqmrE6hpww4g/WcXWY+1hUJ4iZdY9YcWSr53sPj/NrE4R0LX67IFlawOzuuAWkmxkhpb/k
mKuEGLuKXix3llrl+RWf3YFIoqKPDjZkCW7FhA/8hmncC6L4hmWxBoj+hvoROfMFZ4oX7jdpElwz
aojHy45Bikjk6bn8mgI5g2Ze7cZJx8Wa944qw+954MSIwdvY8qBtvaO6A7D6EL1pyezgyTpeI2tl
fqfmQXxMQh9wKwSHDndUm9r6lsL+6iS0FJvbHFTW5G8T8OGan4OxQCbU86QAlccIK2xZzsz116mK
USnbBlc6nwhsOzkqlvy4ec44KE0Uk555dXoOl1O1/JSZ/7yhCyoDQQ5VO8Eqm1EjVg/MTWFMi/Xy
l6ulD4WQpe1SKkT4j9BHZQFFZjqaSrip4p7KqVBs5yI0A4qqqst23vAbLA==
`protect end_protected
